
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"71",x"01",x"01",x"00"),
     1 => (x"00",x"07",x"0f",x"79"),
     2 => (x"49",x"7f",x"36",x"00"),
     3 => (x"00",x"36",x"7f",x"49"),
     4 => (x"49",x"4f",x"06",x"00"),
     5 => (x"00",x"1e",x"3f",x"69"),
     6 => (x"66",x"00",x"00",x"00"),
     7 => (x"00",x"00",x"00",x"66"),
     8 => (x"e6",x"80",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"66"),
    10 => (x"14",x"08",x"08",x"00"),
    11 => (x"00",x"22",x"22",x"14"),
    12 => (x"14",x"14",x"14",x"00"),
    13 => (x"00",x"14",x"14",x"14"),
    14 => (x"14",x"22",x"22",x"00"),
    15 => (x"00",x"08",x"08",x"14"),
    16 => (x"51",x"03",x"02",x"00"),
    17 => (x"00",x"06",x"0f",x"59"),
    18 => (x"5d",x"41",x"7f",x"3e"),
    19 => (x"00",x"1e",x"1f",x"55"),
    20 => (x"09",x"7f",x"7e",x"00"),
    21 => (x"00",x"7e",x"7f",x"09"),
    22 => (x"49",x"7f",x"7f",x"00"),
    23 => (x"00",x"36",x"7f",x"49"),
    24 => (x"63",x"3e",x"1c",x"00"),
    25 => (x"00",x"41",x"41",x"41"),
    26 => (x"41",x"7f",x"7f",x"00"),
    27 => (x"00",x"1c",x"3e",x"63"),
    28 => (x"49",x"7f",x"7f",x"00"),
    29 => (x"00",x"41",x"41",x"49"),
    30 => (x"09",x"7f",x"7f",x"00"),
    31 => (x"00",x"01",x"01",x"09"),
    32 => (x"41",x"7f",x"3e",x"00"),
    33 => (x"00",x"7a",x"7b",x"49"),
    34 => (x"08",x"7f",x"7f",x"00"),
    35 => (x"00",x"7f",x"7f",x"08"),
    36 => (x"7f",x"41",x"00",x"00"),
    37 => (x"00",x"00",x"41",x"7f"),
    38 => (x"40",x"60",x"20",x"00"),
    39 => (x"00",x"3f",x"7f",x"40"),
    40 => (x"1c",x"08",x"7f",x"7f"),
    41 => (x"00",x"41",x"63",x"36"),
    42 => (x"40",x"7f",x"7f",x"00"),
    43 => (x"00",x"40",x"40",x"40"),
    44 => (x"0c",x"06",x"7f",x"7f"),
    45 => (x"00",x"7f",x"7f",x"06"),
    46 => (x"0c",x"06",x"7f",x"7f"),
    47 => (x"00",x"7f",x"7f",x"18"),
    48 => (x"41",x"7f",x"3e",x"00"),
    49 => (x"00",x"3e",x"7f",x"41"),
    50 => (x"09",x"7f",x"7f",x"00"),
    51 => (x"00",x"06",x"0f",x"09"),
    52 => (x"61",x"41",x"7f",x"3e"),
    53 => (x"00",x"40",x"7e",x"7f"),
    54 => (x"09",x"7f",x"7f",x"00"),
    55 => (x"00",x"66",x"7f",x"19"),
    56 => (x"4d",x"6f",x"26",x"00"),
    57 => (x"00",x"32",x"7b",x"59"),
    58 => (x"7f",x"01",x"01",x"00"),
    59 => (x"00",x"01",x"01",x"7f"),
    60 => (x"40",x"7f",x"3f",x"00"),
    61 => (x"00",x"3f",x"7f",x"40"),
    62 => (x"70",x"3f",x"0f",x"00"),
    63 => (x"00",x"0f",x"3f",x"70"),
    64 => (x"18",x"30",x"7f",x"7f"),
    65 => (x"00",x"7f",x"7f",x"30"),
    66 => (x"1c",x"36",x"63",x"41"),
    67 => (x"41",x"63",x"36",x"1c"),
    68 => (x"7c",x"06",x"03",x"01"),
    69 => (x"01",x"03",x"06",x"7c"),
    70 => (x"4d",x"59",x"71",x"61"),
    71 => (x"00",x"41",x"43",x"47"),
    72 => (x"7f",x"7f",x"00",x"00"),
    73 => (x"00",x"00",x"41",x"41"),
    74 => (x"0c",x"06",x"03",x"01"),
    75 => (x"40",x"60",x"30",x"18"),
    76 => (x"41",x"41",x"00",x"00"),
    77 => (x"00",x"00",x"7f",x"7f"),
    78 => (x"03",x"06",x"0c",x"08"),
    79 => (x"00",x"08",x"0c",x"06"),
    80 => (x"80",x"80",x"80",x"80"),
    81 => (x"00",x"80",x"80",x"80"),
    82 => (x"03",x"00",x"00",x"00"),
    83 => (x"00",x"00",x"04",x"07"),
    84 => (x"54",x"74",x"20",x"00"),
    85 => (x"00",x"78",x"7c",x"54"),
    86 => (x"44",x"7f",x"7f",x"00"),
    87 => (x"00",x"38",x"7c",x"44"),
    88 => (x"44",x"7c",x"38",x"00"),
    89 => (x"00",x"00",x"44",x"44"),
    90 => (x"44",x"7c",x"38",x"00"),
    91 => (x"00",x"7f",x"7f",x"44"),
    92 => (x"54",x"7c",x"38",x"00"),
    93 => (x"00",x"18",x"5c",x"54"),
    94 => (x"7f",x"7e",x"04",x"00"),
    95 => (x"00",x"00",x"05",x"05"),
    96 => (x"a4",x"bc",x"18",x"00"),
    97 => (x"00",x"7c",x"fc",x"a4"),
    98 => (x"04",x"7f",x"7f",x"00"),
    99 => (x"00",x"78",x"7c",x"04"),
   100 => (x"3d",x"00",x"00",x"00"),
   101 => (x"00",x"00",x"40",x"7d"),
   102 => (x"80",x"80",x"80",x"00"),
   103 => (x"00",x"00",x"7d",x"fd"),
   104 => (x"10",x"7f",x"7f",x"00"),
   105 => (x"00",x"44",x"6c",x"38"),
   106 => (x"3f",x"00",x"00",x"00"),
   107 => (x"00",x"00",x"40",x"7f"),
   108 => (x"18",x"0c",x"7c",x"7c"),
   109 => (x"00",x"78",x"7c",x"0c"),
   110 => (x"04",x"7c",x"7c",x"00"),
   111 => (x"00",x"78",x"7c",x"04"),
   112 => (x"44",x"7c",x"38",x"00"),
   113 => (x"00",x"38",x"7c",x"44"),
   114 => (x"24",x"fc",x"fc",x"00"),
   115 => (x"00",x"18",x"3c",x"24"),
   116 => (x"24",x"3c",x"18",x"00"),
   117 => (x"00",x"fc",x"fc",x"24"),
   118 => (x"04",x"7c",x"7c",x"00"),
   119 => (x"00",x"08",x"0c",x"04"),
   120 => (x"54",x"5c",x"48",x"00"),
   121 => (x"00",x"20",x"74",x"54"),
   122 => (x"7f",x"3f",x"04",x"00"),
   123 => (x"00",x"00",x"44",x"44"),
   124 => (x"40",x"7c",x"3c",x"00"),
   125 => (x"00",x"7c",x"7c",x"40"),
   126 => (x"60",x"3c",x"1c",x"00"),
   127 => (x"00",x"1c",x"3c",x"60"),
   128 => (x"30",x"60",x"7c",x"3c"),
   129 => (x"00",x"3c",x"7c",x"60"),
   130 => (x"10",x"38",x"6c",x"44"),
   131 => (x"00",x"44",x"6c",x"38"),
   132 => (x"e0",x"bc",x"1c",x"00"),
   133 => (x"00",x"1c",x"3c",x"60"),
   134 => (x"74",x"64",x"44",x"00"),
   135 => (x"00",x"44",x"4c",x"5c"),
   136 => (x"3e",x"08",x"08",x"00"),
   137 => (x"00",x"41",x"41",x"77"),
   138 => (x"7f",x"00",x"00",x"00"),
   139 => (x"00",x"00",x"00",x"7f"),
   140 => (x"77",x"41",x"41",x"00"),
   141 => (x"00",x"08",x"08",x"3e"),
   142 => (x"03",x"01",x"01",x"02"),
   143 => (x"00",x"01",x"02",x"02"),
   144 => (x"7f",x"7f",x"7f",x"7f"),
   145 => (x"00",x"7f",x"7f",x"7f"),
   146 => (x"1c",x"1c",x"08",x"08"),
   147 => (x"7f",x"7f",x"3e",x"3e"),
   148 => (x"3e",x"3e",x"7f",x"7f"),
   149 => (x"08",x"08",x"1c",x"1c"),
   150 => (x"7c",x"18",x"10",x"00"),
   151 => (x"00",x"10",x"18",x"7c"),
   152 => (x"7c",x"30",x"10",x"00"),
   153 => (x"00",x"10",x"30",x"7c"),
   154 => (x"60",x"60",x"30",x"10"),
   155 => (x"00",x"06",x"1e",x"78"),
   156 => (x"18",x"3c",x"66",x"42"),
   157 => (x"00",x"42",x"66",x"3c"),
   158 => (x"c2",x"6a",x"38",x"78"),
   159 => (x"00",x"38",x"6c",x"c6"),
   160 => (x"60",x"00",x"00",x"60"),
   161 => (x"00",x"60",x"00",x"00"),
   162 => (x"5c",x"5b",x"5e",x"0e"),
   163 => (x"86",x"fc",x"0e",x"5d"),
   164 => (x"f2",x"c2",x"7e",x"71"),
   165 => (x"c0",x"4c",x"bf",x"ec"),
   166 => (x"c4",x"1e",x"c0",x"4b"),
   167 => (x"c4",x"02",x"ab",x"66"),
   168 => (x"c2",x"4d",x"c0",x"87"),
   169 => (x"75",x"4d",x"c1",x"87"),
   170 => (x"ee",x"49",x"73",x"1e"),
   171 => (x"86",x"c8",x"87",x"e1"),
   172 => (x"ef",x"49",x"e0",x"c0"),
   173 => (x"a4",x"c4",x"87",x"ea"),
   174 => (x"f0",x"49",x"6a",x"4a"),
   175 => (x"c8",x"f1",x"87",x"f1"),
   176 => (x"c1",x"84",x"cc",x"87"),
   177 => (x"ab",x"b7",x"c8",x"83"),
   178 => (x"87",x"cd",x"ff",x"04"),
   179 => (x"4d",x"26",x"8e",x"fc"),
   180 => (x"4b",x"26",x"4c",x"26"),
   181 => (x"71",x"1e",x"4f",x"26"),
   182 => (x"f0",x"f2",x"c2",x"4a"),
   183 => (x"f0",x"f2",x"c2",x"5a"),
   184 => (x"49",x"78",x"c7",x"48"),
   185 => (x"26",x"87",x"e1",x"fe"),
   186 => (x"1e",x"73",x"1e",x"4f"),
   187 => (x"b7",x"c0",x"4a",x"71"),
   188 => (x"87",x"d3",x"03",x"aa"),
   189 => (x"bf",x"cc",x"d8",x"c2"),
   190 => (x"c1",x"87",x"c4",x"05"),
   191 => (x"c0",x"87",x"c2",x"4b"),
   192 => (x"d0",x"d8",x"c2",x"4b"),
   193 => (x"c2",x"87",x"c4",x"5b"),
   194 => (x"fc",x"5a",x"d0",x"d8"),
   195 => (x"cc",x"d8",x"c2",x"48"),
   196 => (x"c1",x"4a",x"78",x"bf"),
   197 => (x"a2",x"c0",x"c1",x"9a"),
   198 => (x"87",x"e6",x"ec",x"49"),
   199 => (x"4f",x"26",x"4b",x"26"),
   200 => (x"c4",x"4a",x"71",x"1e"),
   201 => (x"49",x"72",x"1e",x"66"),
   202 => (x"fc",x"87",x"f0",x"eb"),
   203 => (x"1e",x"4f",x"26",x"8e"),
   204 => (x"c3",x"48",x"d4",x"ff"),
   205 => (x"d0",x"ff",x"78",x"ff"),
   206 => (x"78",x"e1",x"c0",x"48"),
   207 => (x"c1",x"48",x"d4",x"ff"),
   208 => (x"c4",x"48",x"71",x"78"),
   209 => (x"08",x"d4",x"ff",x"30"),
   210 => (x"48",x"d0",x"ff",x"78"),
   211 => (x"26",x"78",x"e0",x"c0"),
   212 => (x"5b",x"5e",x"0e",x"4f"),
   213 => (x"f0",x"0e",x"5d",x"5c"),
   214 => (x"48",x"a6",x"c8",x"86"),
   215 => (x"ec",x"4d",x"78",x"c0"),
   216 => (x"80",x"fc",x"7e",x"bf"),
   217 => (x"bf",x"ec",x"f2",x"c2"),
   218 => (x"4c",x"bf",x"e8",x"78"),
   219 => (x"bf",x"cc",x"d8",x"c2"),
   220 => (x"87",x"e9",x"e4",x"49"),
   221 => (x"ca",x"49",x"ee",x"cb"),
   222 => (x"4b",x"70",x"87",x"d6"),
   223 => (x"e2",x"e7",x"49",x"c7"),
   224 => (x"05",x"98",x"70",x"87"),
   225 => (x"49",x"6e",x"87",x"c8"),
   226 => (x"c1",x"02",x"99",x"c1"),
   227 => (x"4d",x"c1",x"87",x"c1"),
   228 => (x"c2",x"7e",x"bf",x"ec"),
   229 => (x"49",x"bf",x"cc",x"d8"),
   230 => (x"73",x"87",x"c2",x"e4"),
   231 => (x"87",x"fc",x"c9",x"49"),
   232 => (x"d7",x"02",x"98",x"70"),
   233 => (x"c4",x"d8",x"c2",x"87"),
   234 => (x"b9",x"c1",x"49",x"bf"),
   235 => (x"59",x"c8",x"d8",x"c2"),
   236 => (x"87",x"fb",x"fd",x"71"),
   237 => (x"c9",x"49",x"ee",x"cb"),
   238 => (x"4b",x"70",x"87",x"d6"),
   239 => (x"e2",x"e6",x"49",x"c7"),
   240 => (x"05",x"98",x"70",x"87"),
   241 => (x"6e",x"87",x"c7",x"ff"),
   242 => (x"05",x"99",x"c1",x"49"),
   243 => (x"75",x"87",x"ff",x"fe"),
   244 => (x"e3",x"c0",x"02",x"9d"),
   245 => (x"cc",x"d8",x"c2",x"87"),
   246 => (x"ba",x"c1",x"4a",x"bf"),
   247 => (x"5a",x"d0",x"d8",x"c2"),
   248 => (x"0a",x"7a",x"0a",x"fc"),
   249 => (x"c0",x"c1",x"9a",x"c1"),
   250 => (x"d5",x"e9",x"49",x"a2"),
   251 => (x"49",x"da",x"c1",x"87"),
   252 => (x"c8",x"87",x"f0",x"e5"),
   253 => (x"78",x"c1",x"48",x"a6"),
   254 => (x"bf",x"cc",x"d8",x"c2"),
   255 => (x"87",x"e9",x"c0",x"05"),
   256 => (x"ff",x"c3",x"49",x"74"),
   257 => (x"c0",x"1e",x"71",x"99"),
   258 => (x"87",x"d4",x"fc",x"49"),
   259 => (x"b7",x"c8",x"49",x"74"),
   260 => (x"c1",x"1e",x"71",x"29"),
   261 => (x"87",x"c8",x"fc",x"49"),
   262 => (x"fd",x"c3",x"86",x"c8"),
   263 => (x"87",x"c3",x"e5",x"49"),
   264 => (x"e4",x"49",x"fa",x"c3"),
   265 => (x"d1",x"c7",x"87",x"fd"),
   266 => (x"c3",x"49",x"74",x"87"),
   267 => (x"b7",x"c8",x"99",x"ff"),
   268 => (x"74",x"b4",x"71",x"2c"),
   269 => (x"87",x"df",x"02",x"9c"),
   270 => (x"bf",x"c8",x"d8",x"c2"),
   271 => (x"87",x"dc",x"c7",x"49"),
   272 => (x"c0",x"05",x"98",x"70"),
   273 => (x"4c",x"c0",x"87",x"c4"),
   274 => (x"e0",x"c2",x"87",x"d3"),
   275 => (x"87",x"c0",x"c7",x"49"),
   276 => (x"58",x"cc",x"d8",x"c2"),
   277 => (x"c2",x"87",x"c6",x"c0"),
   278 => (x"c0",x"48",x"c8",x"d8"),
   279 => (x"c8",x"49",x"74",x"78"),
   280 => (x"87",x"ce",x"05",x"99"),
   281 => (x"e3",x"49",x"f5",x"c3"),
   282 => (x"49",x"70",x"87",x"f9"),
   283 => (x"c0",x"02",x"99",x"c2"),
   284 => (x"f2",x"c2",x"87",x"e9"),
   285 => (x"c0",x"02",x"bf",x"f0"),
   286 => (x"c1",x"48",x"87",x"c9"),
   287 => (x"f4",x"f2",x"c2",x"88"),
   288 => (x"c4",x"87",x"d3",x"58"),
   289 => (x"e0",x"c1",x"48",x"66"),
   290 => (x"6e",x"7e",x"70",x"80"),
   291 => (x"c5",x"c0",x"02",x"bf"),
   292 => (x"49",x"ff",x"4b",x"87"),
   293 => (x"a6",x"c8",x"0f",x"73"),
   294 => (x"74",x"78",x"c1",x"48"),
   295 => (x"05",x"99",x"c4",x"49"),
   296 => (x"c3",x"87",x"ce",x"c0"),
   297 => (x"fa",x"e2",x"49",x"f2"),
   298 => (x"c2",x"49",x"70",x"87"),
   299 => (x"f0",x"c0",x"02",x"99"),
   300 => (x"f0",x"f2",x"c2",x"87"),
   301 => (x"c7",x"48",x"7e",x"bf"),
   302 => (x"c0",x"03",x"a8",x"b7"),
   303 => (x"48",x"6e",x"87",x"cb"),
   304 => (x"f2",x"c2",x"80",x"c1"),
   305 => (x"d3",x"c0",x"58",x"f4"),
   306 => (x"48",x"66",x"c4",x"87"),
   307 => (x"70",x"80",x"e0",x"c1"),
   308 => (x"02",x"bf",x"6e",x"7e"),
   309 => (x"4b",x"87",x"c5",x"c0"),
   310 => (x"0f",x"73",x"49",x"fe"),
   311 => (x"c1",x"48",x"a6",x"c8"),
   312 => (x"49",x"fd",x"c3",x"78"),
   313 => (x"70",x"87",x"fc",x"e1"),
   314 => (x"02",x"99",x"c2",x"49"),
   315 => (x"c2",x"87",x"e9",x"c0"),
   316 => (x"02",x"bf",x"f0",x"f2"),
   317 => (x"c2",x"87",x"c9",x"c0"),
   318 => (x"c0",x"48",x"f0",x"f2"),
   319 => (x"87",x"d3",x"c0",x"78"),
   320 => (x"c1",x"48",x"66",x"c4"),
   321 => (x"7e",x"70",x"80",x"e0"),
   322 => (x"c0",x"02",x"bf",x"6e"),
   323 => (x"fd",x"4b",x"87",x"c5"),
   324 => (x"c8",x"0f",x"73",x"49"),
   325 => (x"78",x"c1",x"48",x"a6"),
   326 => (x"e1",x"49",x"fa",x"c3"),
   327 => (x"49",x"70",x"87",x"c5"),
   328 => (x"c0",x"02",x"99",x"c2"),
   329 => (x"f2",x"c2",x"87",x"ea"),
   330 => (x"c7",x"48",x"bf",x"f0"),
   331 => (x"c0",x"03",x"a8",x"b7"),
   332 => (x"f2",x"c2",x"87",x"c9"),
   333 => (x"78",x"c7",x"48",x"f0"),
   334 => (x"c4",x"87",x"d0",x"c0"),
   335 => (x"e0",x"c1",x"4a",x"66"),
   336 => (x"c0",x"02",x"6a",x"82"),
   337 => (x"fc",x"4b",x"87",x"c5"),
   338 => (x"c8",x"0f",x"73",x"49"),
   339 => (x"78",x"c1",x"48",x"a6"),
   340 => (x"f2",x"c2",x"4d",x"c0"),
   341 => (x"50",x"c0",x"48",x"e8"),
   342 => (x"c2",x"49",x"ee",x"cb"),
   343 => (x"4b",x"70",x"87",x"f2"),
   344 => (x"97",x"e8",x"f2",x"c2"),
   345 => (x"dd",x"c1",x"05",x"bf"),
   346 => (x"c3",x"49",x"74",x"87"),
   347 => (x"c0",x"05",x"99",x"f0"),
   348 => (x"da",x"c1",x"87",x"cd"),
   349 => (x"ea",x"df",x"ff",x"49"),
   350 => (x"02",x"98",x"70",x"87"),
   351 => (x"c1",x"87",x"c7",x"c1"),
   352 => (x"4c",x"bf",x"e8",x"4d"),
   353 => (x"99",x"ff",x"c3",x"49"),
   354 => (x"71",x"2c",x"b7",x"c8"),
   355 => (x"cc",x"d8",x"c2",x"b4"),
   356 => (x"dc",x"ff",x"49",x"bf"),
   357 => (x"49",x"73",x"87",x"c7"),
   358 => (x"70",x"87",x"c1",x"c2"),
   359 => (x"c6",x"c0",x"02",x"98"),
   360 => (x"e8",x"f2",x"c2",x"87"),
   361 => (x"c2",x"50",x"c1",x"48"),
   362 => (x"bf",x"97",x"e8",x"f2"),
   363 => (x"87",x"d6",x"c0",x"05"),
   364 => (x"f0",x"c3",x"49",x"74"),
   365 => (x"c6",x"ff",x"05",x"99"),
   366 => (x"49",x"da",x"c1",x"87"),
   367 => (x"87",x"e3",x"de",x"ff"),
   368 => (x"fe",x"05",x"98",x"70"),
   369 => (x"9d",x"75",x"87",x"f9"),
   370 => (x"87",x"e0",x"c0",x"02"),
   371 => (x"c2",x"48",x"a6",x"cc"),
   372 => (x"78",x"bf",x"f0",x"f2"),
   373 => (x"cc",x"49",x"66",x"cc"),
   374 => (x"48",x"66",x"c4",x"91"),
   375 => (x"7e",x"70",x"80",x"71"),
   376 => (x"c0",x"02",x"bf",x"6e"),
   377 => (x"cc",x"4b",x"87",x"c6"),
   378 => (x"0f",x"73",x"49",x"66"),
   379 => (x"c0",x"02",x"66",x"c8"),
   380 => (x"f2",x"c2",x"87",x"c8"),
   381 => (x"f2",x"49",x"bf",x"f0"),
   382 => (x"8e",x"f0",x"87",x"ce"),
   383 => (x"4c",x"26",x"4d",x"26"),
   384 => (x"4f",x"26",x"4b",x"26"),
   385 => (x"00",x"00",x"00",x"00"),
   386 => (x"00",x"00",x"00",x"00"),
   387 => (x"00",x"00",x"00",x"00"),
   388 => (x"ff",x"4a",x"71",x"1e"),
   389 => (x"72",x"49",x"bf",x"c8"),
   390 => (x"4f",x"26",x"48",x"a1"),
   391 => (x"bf",x"c8",x"ff",x"1e"),
   392 => (x"c0",x"c0",x"fe",x"89"),
   393 => (x"a9",x"c0",x"c0",x"c0"),
   394 => (x"c0",x"87",x"c4",x"01"),
   395 => (x"c1",x"87",x"c2",x"4a"),
   396 => (x"26",x"48",x"72",x"4a"),
   397 => (x"5b",x"5e",x"0e",x"4f"),
   398 => (x"71",x"0e",x"5d",x"5c"),
   399 => (x"4c",x"d4",x"ff",x"4b"),
   400 => (x"c0",x"48",x"66",x"d0"),
   401 => (x"ff",x"49",x"d6",x"78"),
   402 => (x"c3",x"87",x"d5",x"de"),
   403 => (x"49",x"6c",x"7c",x"ff"),
   404 => (x"71",x"99",x"ff",x"c3"),
   405 => (x"f0",x"c3",x"49",x"4d"),
   406 => (x"a9",x"e0",x"c1",x"99"),
   407 => (x"c3",x"87",x"cb",x"05"),
   408 => (x"48",x"6c",x"7c",x"ff"),
   409 => (x"66",x"d0",x"98",x"c3"),
   410 => (x"ff",x"c3",x"78",x"08"),
   411 => (x"49",x"4a",x"6c",x"7c"),
   412 => (x"ff",x"c3",x"31",x"c8"),
   413 => (x"71",x"4a",x"6c",x"7c"),
   414 => (x"c8",x"49",x"72",x"b2"),
   415 => (x"7c",x"ff",x"c3",x"31"),
   416 => (x"b2",x"71",x"4a",x"6c"),
   417 => (x"31",x"c8",x"49",x"72"),
   418 => (x"6c",x"7c",x"ff",x"c3"),
   419 => (x"ff",x"b2",x"71",x"4a"),
   420 => (x"e0",x"c0",x"48",x"d0"),
   421 => (x"02",x"9b",x"73",x"78"),
   422 => (x"7b",x"72",x"87",x"c2"),
   423 => (x"4d",x"26",x"48",x"75"),
   424 => (x"4b",x"26",x"4c",x"26"),
   425 => (x"26",x"1e",x"4f",x"26"),
   426 => (x"5b",x"5e",x"0e",x"4f"),
   427 => (x"86",x"f8",x"0e",x"5c"),
   428 => (x"a6",x"c8",x"1e",x"76"),
   429 => (x"87",x"fd",x"fd",x"49"),
   430 => (x"4b",x"70",x"86",x"c4"),
   431 => (x"a8",x"c2",x"48",x"6e"),
   432 => (x"87",x"f0",x"c2",x"03"),
   433 => (x"f0",x"c3",x"4a",x"73"),
   434 => (x"aa",x"d0",x"c1",x"9a"),
   435 => (x"c1",x"87",x"c7",x"02"),
   436 => (x"c2",x"05",x"aa",x"e0"),
   437 => (x"49",x"73",x"87",x"de"),
   438 => (x"c3",x"02",x"99",x"c8"),
   439 => (x"87",x"c6",x"ff",x"87"),
   440 => (x"9c",x"c3",x"4c",x"73"),
   441 => (x"c1",x"05",x"ac",x"c2"),
   442 => (x"66",x"c4",x"87",x"c2"),
   443 => (x"71",x"31",x"c9",x"49"),
   444 => (x"4a",x"66",x"c4",x"1e"),
   445 => (x"f2",x"c2",x"92",x"d4"),
   446 => (x"81",x"72",x"49",x"f4"),
   447 => (x"87",x"d9",x"cf",x"fe"),
   448 => (x"db",x"ff",x"49",x"d8"),
   449 => (x"c0",x"c8",x"87",x"da"),
   450 => (x"cc",x"e1",x"c2",x"1e"),
   451 => (x"c6",x"e9",x"fd",x"49"),
   452 => (x"48",x"d0",x"ff",x"87"),
   453 => (x"c2",x"78",x"e0",x"c0"),
   454 => (x"cc",x"1e",x"cc",x"e1"),
   455 => (x"92",x"d4",x"4a",x"66"),
   456 => (x"49",x"f4",x"f2",x"c2"),
   457 => (x"cd",x"fe",x"81",x"72"),
   458 => (x"86",x"cc",x"87",x"e0"),
   459 => (x"c1",x"05",x"ac",x"c1"),
   460 => (x"66",x"c4",x"87",x"c2"),
   461 => (x"71",x"31",x"c9",x"49"),
   462 => (x"4a",x"66",x"c4",x"1e"),
   463 => (x"f2",x"c2",x"92",x"d4"),
   464 => (x"81",x"72",x"49",x"f4"),
   465 => (x"87",x"d1",x"ce",x"fe"),
   466 => (x"1e",x"cc",x"e1",x"c2"),
   467 => (x"d4",x"4a",x"66",x"c8"),
   468 => (x"f4",x"f2",x"c2",x"92"),
   469 => (x"fe",x"81",x"72",x"49"),
   470 => (x"d7",x"87",x"e0",x"cb"),
   471 => (x"ff",x"d9",x"ff",x"49"),
   472 => (x"1e",x"c0",x"c8",x"87"),
   473 => (x"49",x"cc",x"e1",x"c2"),
   474 => (x"87",x"c8",x"e7",x"fd"),
   475 => (x"d0",x"ff",x"86",x"cc"),
   476 => (x"78",x"e0",x"c0",x"48"),
   477 => (x"4c",x"26",x"8e",x"f8"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"86",x"fc",x"0e",x"5d"),
   481 => (x"d4",x"ff",x"4d",x"71"),
   482 => (x"7e",x"66",x"d4",x"4c"),
   483 => (x"a8",x"b7",x"c3",x"48"),
   484 => (x"87",x"e2",x"c1",x"01"),
   485 => (x"66",x"c4",x"1e",x"75"),
   486 => (x"c2",x"93",x"d4",x"4b"),
   487 => (x"73",x"83",x"f4",x"f2"),
   488 => (x"d0",x"c5",x"fe",x"49"),
   489 => (x"49",x"a3",x"c8",x"87"),
   490 => (x"d0",x"ff",x"49",x"69"),
   491 => (x"78",x"e1",x"c8",x"48"),
   492 => (x"48",x"71",x"7c",x"dd"),
   493 => (x"70",x"98",x"ff",x"c3"),
   494 => (x"c8",x"4a",x"71",x"7c"),
   495 => (x"48",x"72",x"2a",x"b7"),
   496 => (x"70",x"98",x"ff",x"c3"),
   497 => (x"d0",x"4a",x"71",x"7c"),
   498 => (x"48",x"72",x"2a",x"b7"),
   499 => (x"70",x"98",x"ff",x"c3"),
   500 => (x"d8",x"48",x"71",x"7c"),
   501 => (x"7c",x"70",x"28",x"b7"),
   502 => (x"7c",x"7c",x"7c",x"c0"),
   503 => (x"7c",x"7c",x"7c",x"7c"),
   504 => (x"7c",x"7c",x"7c",x"7c"),
   505 => (x"48",x"d0",x"ff",x"7c"),
   506 => (x"c4",x"78",x"e0",x"c0"),
   507 => (x"49",x"dc",x"1e",x"66"),
   508 => (x"87",x"d1",x"d8",x"ff"),
   509 => (x"8e",x"fc",x"86",x"c8"),
   510 => (x"4c",x"26",x"4d",x"26"),
   511 => (x"4f",x"26",x"4b",x"26"),
   512 => (x"d0",x"e0",x"c2",x"1e"),
   513 => (x"de",x"fe",x"49",x"bf"),
   514 => (x"48",x"c0",x"87",x"c0"),
   515 => (x"00",x"00",x"4f",x"26"),
   516 => (x"00",x"00",x"28",x"14"),
   517 => (x"32",x"43",x"49",x"56"),
   518 => (x"20",x"20",x"20",x"30"),
   519 => (x"00",x"4d",x"4f",x"52"),
   520 => (x"00",x"00",x"1b",x"b3"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

