library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dcf3c287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49dcf3c2",
    18 => x"48e4e0c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"e4e0c287",
    25 => x"e0e0c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e8c187f7",
    29 => x"e0c287ca",
    30 => x"e0c24de4",
    31 => x"ad744ce4",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"711e731e",
    78 => x"4b66c84a",
    79 => x"718bc149",
    80 => x"87cf0299",
    81 => x"d4ff4812",
    82 => x"49737808",
    83 => x"99718bc1",
    84 => x"2687f105",
    85 => x"0e4f264b",
    86 => x"0e5c5b5e",
    87 => x"d4ff4a71",
    88 => x"4b66cc4c",
    89 => x"718bc149",
    90 => x"87ce0299",
    91 => x"6c7cffc3",
    92 => x"c1497352",
    93 => x"0599718b",
    94 => x"4c2687f2",
    95 => x"4f264b26",
    96 => x"ff1e731e",
    97 => x"ffc34bd4",
    98 => x"c34a6b7b",
    99 => x"496b7bff",
   100 => x"b17232c8",
   101 => x"6b7bffc3",
   102 => x"7131c84a",
   103 => x"7bffc3b2",
   104 => x"32c8496b",
   105 => x"4871b172",
   106 => x"4f264b26",
   107 => x"5c5b5e0e",
   108 => x"4d710e5d",
   109 => x"754cd4ff",
   110 => x"98ffc348",
   111 => x"e0c27c70",
   112 => x"c805bfe4",
   113 => x"4866d087",
   114 => x"a6d430c9",
   115 => x"4966d058",
   116 => x"487129d8",
   117 => x"7098ffc3",
   118 => x"4966d07c",
   119 => x"487129d0",
   120 => x"7098ffc3",
   121 => x"4966d07c",
   122 => x"487129c8",
   123 => x"7098ffc3",
   124 => x"4866d07c",
   125 => x"7098ffc3",
   126 => x"d049757c",
   127 => x"c3487129",
   128 => x"7c7098ff",
   129 => x"f0c94b6c",
   130 => x"ffc34aff",
   131 => x"87cf05ab",
   132 => x"6c7c7149",
   133 => x"028ac14b",
   134 => x"ab7187c5",
   135 => x"7387f202",
   136 => x"264d2648",
   137 => x"264b264c",
   138 => x"49c01e4f",
   139 => x"c348d4ff",
   140 => x"81c178ff",
   141 => x"a9b7c8c3",
   142 => x"2687f104",
   143 => x"5b5e0e4f",
   144 => x"c00e5d5c",
   145 => x"f7c1f0ff",
   146 => x"c0c0c14d",
   147 => x"4bc0c0c0",
   148 => x"c487d6ff",
   149 => x"c04cdff8",
   150 => x"fd49751e",
   151 => x"86c487ce",
   152 => x"c005a8c1",
   153 => x"d4ff87e5",
   154 => x"78ffc348",
   155 => x"e1c01e73",
   156 => x"49e9c1f0",
   157 => x"c487f5fc",
   158 => x"05987086",
   159 => x"d4ff87ca",
   160 => x"78ffc348",
   161 => x"87cb48c1",
   162 => x"c187defe",
   163 => x"c6ff058c",
   164 => x"2648c087",
   165 => x"264c264d",
   166 => x"0e4f264b",
   167 => x"0e5c5b5e",
   168 => x"c1f0ffc0",
   169 => x"d4ff4cc1",
   170 => x"78ffc348",
   171 => x"f749e0cb",
   172 => x"4bd387f5",
   173 => x"49741ec0",
   174 => x"c487f1fb",
   175 => x"05987086",
   176 => x"d4ff87ca",
   177 => x"78ffc348",
   178 => x"87cb48c1",
   179 => x"c187dafd",
   180 => x"dfff058b",
   181 => x"2648c087",
   182 => x"264b264c",
   183 => x"0000004f",
   184 => x"00444d43",
   185 => x"5c5b5e0e",
   186 => x"ffc30e5d",
   187 => x"4bd4ff4d",
   188 => x"c687f6fc",
   189 => x"e1c01eea",
   190 => x"49c8c1f0",
   191 => x"c487edfa",
   192 => x"02a8c186",
   193 => x"d2fe87c8",
   194 => x"c148c087",
   195 => x"eff987e8",
   196 => x"cf497087",
   197 => x"c699ffff",
   198 => x"c802a9ea",
   199 => x"87fbfd87",
   200 => x"d1c148c0",
   201 => x"c07b7587",
   202 => x"d0fc4cf1",
   203 => x"02987087",
   204 => x"c087ecc0",
   205 => x"f0ffc01e",
   206 => x"f949fac1",
   207 => x"86c487ee",
   208 => x"da059870",
   209 => x"6b7b7587",
   210 => x"757b7549",
   211 => x"757b757b",
   212 => x"99c0c17b",
   213 => x"c187c402",
   214 => x"c087db48",
   215 => x"c287d748",
   216 => x"87ca05ac",
   217 => x"f449c0ce",
   218 => x"48c087fd",
   219 => x"8cc187c8",
   220 => x"87f6fe05",
   221 => x"4d2648c0",
   222 => x"4b264c26",
   223 => x"00004f26",
   224 => x"43484453",
   225 => x"69616620",
   226 => x"000a216c",
   227 => x"5c5b5e0e",
   228 => x"d0ff0e5d",
   229 => x"d0e5c04d",
   230 => x"c24cc0c1",
   231 => x"c148e4e0",
   232 => x"49d8d078",
   233 => x"c787c0f4",
   234 => x"f97dc24b",
   235 => x"7dc387fb",
   236 => x"49741ec0",
   237 => x"c487f5f7",
   238 => x"05a8c186",
   239 => x"c24b87c1",
   240 => x"87cb05ab",
   241 => x"f349d0d0",
   242 => x"48c087dd",
   243 => x"c187f6c0",
   244 => x"d4ff058b",
   245 => x"87ccfc87",
   246 => x"58e8e0c2",
   247 => x"cd059870",
   248 => x"c01ec187",
   249 => x"d0c1f0ff",
   250 => x"87c0f749",
   251 => x"d4ff86c4",
   252 => x"78ffc348",
   253 => x"c287ccc5",
   254 => x"c258ece0",
   255 => x"48d4ff7d",
   256 => x"c178ffc3",
   257 => x"264d2648",
   258 => x"264b264c",
   259 => x"0000004f",
   260 => x"52524549",
   261 => x"00000000",
   262 => x"00495053",
   263 => x"5c5b5e0e",
   264 => x"4d710e5d",
   265 => x"ff4cffc3",
   266 => x"7b744bd4",
   267 => x"c448d0ff",
   268 => x"7b7478c3",
   269 => x"ffc01e75",
   270 => x"49d8c1f0",
   271 => x"c487edf5",
   272 => x"02987086",
   273 => x"c8d287cb",
   274 => x"87dbf149",
   275 => x"eec048c1",
   276 => x"c37b7487",
   277 => x"c0c87bfe",
   278 => x"4966d41e",
   279 => x"c487d5f3",
   280 => x"747b7486",
   281 => x"d87b747b",
   282 => x"744ae0da",
   283 => x"c5056b7b",
   284 => x"058ac187",
   285 => x"7b7487f5",
   286 => x"c248d0ff",
   287 => x"2648c078",
   288 => x"264c264d",
   289 => x"004f264b",
   290 => x"74697257",
   291 => x"61662065",
   292 => x"64656c69",
   293 => x"5e0e000a",
   294 => x"0e5d5c5b",
   295 => x"4b7186fc",
   296 => x"c04cd4ff",
   297 => x"cdeec57e",
   298 => x"ffc34adf",
   299 => x"c3486c7c",
   300 => x"c005a8fe",
   301 => x"4d7487f8",
   302 => x"cc029b73",
   303 => x"1e66d487",
   304 => x"d2f24973",
   305 => x"d486c487",
   306 => x"48d0ff87",
   307 => x"d478d1c4",
   308 => x"ffc34a66",
   309 => x"058ac17d",
   310 => x"a6d887f8",
   311 => x"7cffc35a",
   312 => x"059b737c",
   313 => x"d0ff87c5",
   314 => x"c178d048",
   315 => x"8ac17e4a",
   316 => x"87f6fe05",
   317 => x"8efc486e",
   318 => x"4c264d26",
   319 => x"4f264b26",
   320 => x"711e731e",
   321 => x"ff4bc04a",
   322 => x"ffc348d4",
   323 => x"48d0ff78",
   324 => x"ff78c3c4",
   325 => x"ffc348d4",
   326 => x"c01e7278",
   327 => x"d1c1f0ff",
   328 => x"87c8f249",
   329 => x"987086c4",
   330 => x"c887d205",
   331 => x"66cc1ec0",
   332 => x"87e2fd49",
   333 => x"4b7086c4",
   334 => x"c248d0ff",
   335 => x"26487378",
   336 => x"0e4f264b",
   337 => x"5d5c5b5e",
   338 => x"c01ec00e",
   339 => x"c9c1f0ff",
   340 => x"87d8f149",
   341 => x"e0c21ed2",
   342 => x"f9fc49ec",
   343 => x"c086c887",
   344 => x"d284c14c",
   345 => x"f804acb7",
   346 => x"ece0c287",
   347 => x"c349bf97",
   348 => x"c0c199c0",
   349 => x"e7c005a9",
   350 => x"f3e0c287",
   351 => x"d049bf97",
   352 => x"f4e0c231",
   353 => x"c84abf97",
   354 => x"c2b17232",
   355 => x"bf97f5e0",
   356 => x"4c71b14a",
   357 => x"ffffffcf",
   358 => x"ca84c19c",
   359 => x"87e7c134",
   360 => x"97f5e0c2",
   361 => x"31c149bf",
   362 => x"e0c299c6",
   363 => x"4abf97f6",
   364 => x"722ab7c7",
   365 => x"f1e0c2b1",
   366 => x"4d4abf97",
   367 => x"e0c29dcf",
   368 => x"4abf97f2",
   369 => x"32ca9ac3",
   370 => x"97f3e0c2",
   371 => x"33c24bbf",
   372 => x"e0c2b273",
   373 => x"4bbf97f4",
   374 => x"c69bc0c3",
   375 => x"b2732bb7",
   376 => x"48c181c2",
   377 => x"49703071",
   378 => x"307548c1",
   379 => x"4c724d70",
   380 => x"947184c1",
   381 => x"adb7c0c8",
   382 => x"c187cc06",
   383 => x"c82db734",
   384 => x"01adb7c0",
   385 => x"7487f4ff",
   386 => x"264d2648",
   387 => x"264b264c",
   388 => x"5b5e0e4f",
   389 => x"f80e5d5c",
   390 => x"d4e9c286",
   391 => x"c278c048",
   392 => x"c01ecce1",
   393 => x"87d8fb49",
   394 => x"987086c4",
   395 => x"c087c505",
   396 => x"87c0c948",
   397 => x"7ec14dc0",
   398 => x"bfdcf7c0",
   399 => x"c2e2c249",
   400 => x"4bc8714a",
   401 => x"7087dfea",
   402 => x"87c20598",
   403 => x"f7c07ec0",
   404 => x"c249bfd8",
   405 => x"714adee2",
   406 => x"c9ea4bc8",
   407 => x"05987087",
   408 => x"7ec087c2",
   409 => x"fdc0026e",
   410 => x"d2e8c287",
   411 => x"e9c24dbf",
   412 => x"7ebf9fca",
   413 => x"ead6c548",
   414 => x"87c705a8",
   415 => x"bfd2e8c2",
   416 => x"6e87ce4d",
   417 => x"d5e9ca48",
   418 => x"87c502a8",
   419 => x"e3c748c0",
   420 => x"cce1c287",
   421 => x"f949751e",
   422 => x"86c487e6",
   423 => x"c5059870",
   424 => x"c748c087",
   425 => x"f7c087ce",
   426 => x"c249bfd8",
   427 => x"714adee2",
   428 => x"f1e84bc8",
   429 => x"05987087",
   430 => x"e9c287c8",
   431 => x"78c148d4",
   432 => x"f7c087da",
   433 => x"c249bfdc",
   434 => x"714ac2e2",
   435 => x"d5e84bc8",
   436 => x"02987087",
   437 => x"c087c5c0",
   438 => x"87d8c648",
   439 => x"97cae9c2",
   440 => x"d5c149bf",
   441 => x"cdc005a9",
   442 => x"cbe9c287",
   443 => x"c249bf97",
   444 => x"c002a9ea",
   445 => x"48c087c5",
   446 => x"c287f9c5",
   447 => x"bf97cce1",
   448 => x"e9c3487e",
   449 => x"cec002a8",
   450 => x"c3486e87",
   451 => x"c002a8eb",
   452 => x"48c087c5",
   453 => x"c287ddc5",
   454 => x"bf97d7e1",
   455 => x"c0059949",
   456 => x"e1c287cc",
   457 => x"49bf97d8",
   458 => x"c002a9c2",
   459 => x"48c087c5",
   460 => x"c287c1c5",
   461 => x"bf97d9e1",
   462 => x"d0e9c248",
   463 => x"484c7058",
   464 => x"e9c288c1",
   465 => x"e1c258d4",
   466 => x"49bf97da",
   467 => x"e1c28175",
   468 => x"4abf97db",
   469 => x"a17232c8",
   470 => x"e4edc27e",
   471 => x"c2786e48",
   472 => x"bf97dce1",
   473 => x"58a6c848",
   474 => x"bfd4e9c2",
   475 => x"87cfc202",
   476 => x"bfd8f7c0",
   477 => x"dee2c249",
   478 => x"4bc8714a",
   479 => x"7087e7e5",
   480 => x"c5c00298",
   481 => x"c348c087",
   482 => x"e9c287ea",
   483 => x"c24cbfcc",
   484 => x"c25cf8ed",
   485 => x"bf97f1e1",
   486 => x"c231c849",
   487 => x"bf97f0e1",
   488 => x"c249a14a",
   489 => x"bf97f2e1",
   490 => x"7232d04a",
   491 => x"e1c249a1",
   492 => x"4abf97f3",
   493 => x"a17232d8",
   494 => x"9166c449",
   495 => x"bfe4edc2",
   496 => x"ecedc281",
   497 => x"f9e1c259",
   498 => x"c84abf97",
   499 => x"f8e1c232",
   500 => x"a24bbf97",
   501 => x"fae1c24a",
   502 => x"d04bbf97",
   503 => x"4aa27333",
   504 => x"97fbe1c2",
   505 => x"9bcf4bbf",
   506 => x"a27333d8",
   507 => x"f0edc24a",
   508 => x"748ac25a",
   509 => x"f0edc292",
   510 => x"78a17248",
   511 => x"c287c1c1",
   512 => x"bf97dee1",
   513 => x"c231c849",
   514 => x"bf97dde1",
   515 => x"c549a14a",
   516 => x"81ffc731",
   517 => x"edc229c9",
   518 => x"e1c259f8",
   519 => x"4abf97e3",
   520 => x"e1c232c8",
   521 => x"4bbf97e2",
   522 => x"66c44aa2",
   523 => x"c2826e92",
   524 => x"c25af4ed",
   525 => x"c048eced",
   526 => x"e8edc278",
   527 => x"78a17248",
   528 => x"48f8edc2",
   529 => x"bfecedc2",
   530 => x"fcedc278",
   531 => x"f0edc248",
   532 => x"e9c278bf",
   533 => x"c002bfd4",
   534 => x"487487c9",
   535 => x"7e7030c4",
   536 => x"c287c9c0",
   537 => x"48bff4ed",
   538 => x"7e7030c4",
   539 => x"48d8e9c2",
   540 => x"48c1786e",
   541 => x"4d268ef8",
   542 => x"4b264c26",
   543 => x"5e0e4f26",
   544 => x"0e5d5c5b",
   545 => x"e9c24a71",
   546 => x"cb02bfd4",
   547 => x"c74b7287",
   548 => x"c14d722b",
   549 => x"87c99dff",
   550 => x"2bc84b72",
   551 => x"ffc34d72",
   552 => x"e4edc29d",
   553 => x"f7c083bf",
   554 => x"02abbfd4",
   555 => x"f7c087d9",
   556 => x"e1c25bd8",
   557 => x"49731ecc",
   558 => x"c487c5f1",
   559 => x"05987086",
   560 => x"48c087c5",
   561 => x"c287e6c0",
   562 => x"02bfd4e9",
   563 => x"497587d2",
   564 => x"e1c291c4",
   565 => x"4c6981cc",
   566 => x"ffffffcf",
   567 => x"87cb9cff",
   568 => x"91c24975",
   569 => x"81cce1c2",
   570 => x"744c699f",
   571 => x"264d2648",
   572 => x"264b264c",
   573 => x"5b5e0e4f",
   574 => x"f40e5d5c",
   575 => x"59a6cc86",
   576 => x"c50566c8",
   577 => x"c348c087",
   578 => x"66c887c8",
   579 => x"7080c848",
   580 => x"78c0487e",
   581 => x"c70266dc",
   582 => x"9766dc87",
   583 => x"87c505bf",
   584 => x"edc248c0",
   585 => x"c11ec087",
   586 => x"eeca4949",
   587 => x"7086c487",
   588 => x"c0029c4c",
   589 => x"e9c287fc",
   590 => x"66dc4adc",
   591 => x"cadeff49",
   592 => x"02987087",
   593 => x"7487ebc0",
   594 => x"4966dc4a",
   595 => x"deff4bcb",
   596 => x"987087ee",
   597 => x"c087db02",
   598 => x"029c741e",
   599 => x"4dc087c4",
   600 => x"4dc187c2",
   601 => x"f2c94975",
   602 => x"7086c487",
   603 => x"ff059c4c",
   604 => x"9c7487c4",
   605 => x"87d8c102",
   606 => x"6e49a4dc",
   607 => x"da786948",
   608 => x"66c849a4",
   609 => x"c880c448",
   610 => x"699f58a6",
   611 => x"0866c448",
   612 => x"d4e9c278",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"c448496e",
   620 => x"c480bf66",
   621 => x"c8780866",
   622 => x"78c04866",
   623 => x"cc4966c8",
   624 => x"bf66c481",
   625 => x"4966c879",
   626 => x"79c081d0",
   627 => x"87c248c1",
   628 => x"8ef448c0",
   629 => x"4c264d26",
   630 => x"4f264b26",
   631 => x"5c5b5e0e",
   632 => x"4c710e5d",
   633 => x"744d66d0",
   634 => x"c6c1029c",
   635 => x"49a4c887",
   636 => x"fec00269",
   637 => x"6c4a7587",
   638 => x"4da17249",
   639 => x"d0e9c2b9",
   640 => x"baff4abf",
   641 => x"99719972",
   642 => x"87e5c002",
   643 => x"6b4ba4c4",
   644 => x"87eaf949",
   645 => x"e9c27b70",
   646 => x"6c49bfcc",
   647 => x"757c7181",
   648 => x"e9c2b94a",
   649 => x"ff4abfd0",
   650 => x"719972ba",
   651 => x"dbff0599",
   652 => x"267c7587",
   653 => x"264c264d",
   654 => x"1e4f264b",
   655 => x"4b711e73",
   656 => x"87c7029b",
   657 => x"6949a3c8",
   658 => x"c087c505",
   659 => x"87f6c048",
   660 => x"bfe8edc2",
   661 => x"4aa3c449",
   662 => x"8ac24a6a",
   663 => x"bfcce9c2",
   664 => x"49a17292",
   665 => x"bfd0e9c2",
   666 => x"729a6b4a",
   667 => x"f7c049a1",
   668 => x"66c859d8",
   669 => x"c7ea711e",
   670 => x"7086c487",
   671 => x"87c40598",
   672 => x"87c248c0",
   673 => x"4b2648c1",
   674 => x"731e4f26",
   675 => x"9b4b711e",
   676 => x"c887c702",
   677 => x"056949a3",
   678 => x"48c087c5",
   679 => x"c287f6c0",
   680 => x"49bfe8ed",
   681 => x"6a4aa3c4",
   682 => x"c28ac24a",
   683 => x"92bfcce9",
   684 => x"c249a172",
   685 => x"4abfd0e9",
   686 => x"a1729a6b",
   687 => x"d8f7c049",
   688 => x"1e66c859",
   689 => x"87d4e571",
   690 => x"987086c4",
   691 => x"c087c405",
   692 => x"c187c248",
   693 => x"264b2648",
   694 => x"5b5e0e4f",
   695 => x"fc0e5d5c",
   696 => x"d44b7186",
   697 => x"9b734d66",
   698 => x"87ccc102",
   699 => x"6949a3c8",
   700 => x"87c4c102",
   701 => x"c24ca3d0",
   702 => x"49bfd0e9",
   703 => x"4a6cb9ff",
   704 => x"66d47e99",
   705 => x"87cd06a9",
   706 => x"cc7c7bc0",
   707 => x"a3c44aa3",
   708 => x"ca796a49",
   709 => x"f8497287",
   710 => x"66d499c0",
   711 => x"758d714d",
   712 => x"7129c949",
   713 => x"fa49731e",
   714 => x"e1c287f2",
   715 => x"49731ecc",
   716 => x"c887c8fc",
   717 => x"7c66d486",
   718 => x"4d268efc",
   719 => x"4b264c26",
   720 => x"731e4f26",
   721 => x"9b4b711e",
   722 => x"87e4c002",
   723 => x"5bfcedc2",
   724 => x"8ac24a73",
   725 => x"bfcce9c2",
   726 => x"edc29249",
   727 => x"7248bfe8",
   728 => x"c0eec280",
   729 => x"c4487158",
   730 => x"dce9c230",
   731 => x"87edc058",
   732 => x"48f8edc2",
   733 => x"bfecedc2",
   734 => x"fcedc278",
   735 => x"f0edc248",
   736 => x"e9c278bf",
   737 => x"c902bfd4",
   738 => x"cce9c287",
   739 => x"31c449bf",
   740 => x"edc287c7",
   741 => x"c449bff4",
   742 => x"dce9c231",
   743 => x"264b2659",
   744 => x"5b5e0e4f",
   745 => x"4a710e5c",
   746 => x"9a724bc0",
   747 => x"87e0c002",
   748 => x"9f49a2da",
   749 => x"e9c24b69",
   750 => x"cf02bfd4",
   751 => x"49a2d487",
   752 => x"4c49699f",
   753 => x"9cffffc0",
   754 => x"87c234d0",
   755 => x"b3744cc0",
   756 => x"edfd4973",
   757 => x"264c2687",
   758 => x"0e4f264b",
   759 => x"5d5c5b5e",
   760 => x"c886f00e",
   761 => x"ffcf59a6",
   762 => x"4cf8ffff",
   763 => x"66c47ec0",
   764 => x"c287d802",
   765 => x"c048c8e1",
   766 => x"c0e1c278",
   767 => x"fcedc248",
   768 => x"e1c278bf",
   769 => x"edc248c4",
   770 => x"c278bff8",
   771 => x"c048e9e9",
   772 => x"d8e9c250",
   773 => x"e1c249bf",
   774 => x"714abfc8",
   775 => x"cbc403aa",
   776 => x"cf497287",
   777 => x"e9c00599",
   778 => x"d4f7c087",
   779 => x"c0e1c248",
   780 => x"e1c278bf",
   781 => x"e1c21ecc",
   782 => x"c249bfc0",
   783 => x"c148c0e1",
   784 => x"e27178a1",
   785 => x"86c487fa",
   786 => x"48d0f7c0",
   787 => x"78cce1c2",
   788 => x"f7c087cc",
   789 => x"c048bfd0",
   790 => x"f7c080e0",
   791 => x"e1c258d4",
   792 => x"c148bfc8",
   793 => x"cce1c280",
   794 => x"0dd02758",
   795 => x"97bf0000",
   796 => x"029d4dbf",
   797 => x"c387e5c2",
   798 => x"c202ade5",
   799 => x"f7c087de",
   800 => x"cb4bbfd0",
   801 => x"4c1149a3",
   802 => x"c105accf",
   803 => x"497587d2",
   804 => x"89c199df",
   805 => x"e9c291cd",
   806 => x"a3c181dc",
   807 => x"c351124a",
   808 => x"51124aa3",
   809 => x"124aa3c5",
   810 => x"4aa3c751",
   811 => x"a3c95112",
   812 => x"ce51124a",
   813 => x"51124aa3",
   814 => x"124aa3d0",
   815 => x"4aa3d251",
   816 => x"a3d45112",
   817 => x"d651124a",
   818 => x"51124aa3",
   819 => x"124aa3d8",
   820 => x"4aa3dc51",
   821 => x"a3de5112",
   822 => x"c151124a",
   823 => x"87fcc07e",
   824 => x"99c84974",
   825 => x"87edc005",
   826 => x"99d04974",
   827 => x"c087d305",
   828 => x"c00266e0",
   829 => x"497387cc",
   830 => x"0f66e0c0",
   831 => x"c0029870",
   832 => x"056e87d3",
   833 => x"c287c6c0",
   834 => x"c048dce9",
   835 => x"d0f7c050",
   836 => x"ebc248bf",
   837 => x"e9e9c287",
   838 => x"7e50c048",
   839 => x"bfd8e9c2",
   840 => x"c8e1c249",
   841 => x"aa714abf",
   842 => x"87f5fb04",
   843 => x"ffffffcf",
   844 => x"edc24cf8",
   845 => x"c005bffc",
   846 => x"e9c287c8",
   847 => x"c102bfd4",
   848 => x"e1c287fc",
   849 => x"ec49bfc4",
   850 => x"e1c287f4",
   851 => x"a6c458c8",
   852 => x"c4e1c248",
   853 => x"e9c278bf",
   854 => x"c002bfd4",
   855 => x"66c487db",
   856 => x"74997449",
   857 => x"c8c002a9",
   858 => x"48a6c887",
   859 => x"e7c078c0",
   860 => x"48a6c887",
   861 => x"dfc078c1",
   862 => x"4966c487",
   863 => x"99f8ffcf",
   864 => x"c8c002a9",
   865 => x"48a6cc87",
   866 => x"c5c078c0",
   867 => x"48a6cc87",
   868 => x"a6c878c1",
   869 => x"7866cc48",
   870 => x"c00566c8",
   871 => x"66c487e0",
   872 => x"c289c249",
   873 => x"4abfcce9",
   874 => x"e8edc291",
   875 => x"e1c24abf",
   876 => x"a17248c0",
   877 => x"c8e1c278",
   878 => x"f978c048",
   879 => x"48c087d3",
   880 => x"ffffffcf",
   881 => x"8ef04cf8",
   882 => x"4c264d26",
   883 => x"4f264b26",
   884 => x"00000000",
   885 => x"ffffffff",
   886 => x"00000de0",
   887 => x"00000dec",
   888 => x"33544146",
   889 => x"20202032",
   890 => x"00000000",
   891 => x"31544146",
   892 => x"20202036",
   893 => x"d4ff1e00",
   894 => x"78ffc348",
   895 => x"4f264868",
   896 => x"48d4ff1e",
   897 => x"ff78ffc3",
   898 => x"e1c048d0",
   899 => x"48d4ff78",
   900 => x"4f2678d4",
   901 => x"48d0ff1e",
   902 => x"2678e0c0",
   903 => x"d4ff1e4f",
   904 => x"99497087",
   905 => x"c087c602",
   906 => x"f105a9fb",
   907 => x"26487187",
   908 => x"5b5e0e4f",
   909 => x"4b710e5c",
   910 => x"f8fe4cc0",
   911 => x"99497087",
   912 => x"87f9c002",
   913 => x"02a9ecc0",
   914 => x"c087f2c0",
   915 => x"c002a9fb",
   916 => x"66cc87eb",
   917 => x"c703acb7",
   918 => x"0266d087",
   919 => x"537187c2",
   920 => x"c2029971",
   921 => x"fe84c187",
   922 => x"497087cb",
   923 => x"87cd0299",
   924 => x"02a9ecc0",
   925 => x"fbc087c7",
   926 => x"d5ff05a9",
   927 => x"0266d087",
   928 => x"97c087c3",
   929 => x"a9ecc07b",
   930 => x"7487c405",
   931 => x"7487c54a",
   932 => x"8a0ac04a",
   933 => x"4c264872",
   934 => x"4f264b26",
   935 => x"87d5fd1e",
   936 => x"c04a4970",
   937 => x"c904aaf0",
   938 => x"aaf9c087",
   939 => x"c087c301",
   940 => x"c1c18af0",
   941 => x"87c904aa",
   942 => x"01aadac1",
   943 => x"f7c087c3",
   944 => x"2648728a",
   945 => x"5b5e0e4f",
   946 => x"f80e5d5c",
   947 => x"c04c7186",
   948 => x"87ecfc7e",
   949 => x"fdc04bc0",
   950 => x"49bf97e4",
   951 => x"cf04a9c0",
   952 => x"87f9fc87",
   953 => x"fdc083c1",
   954 => x"49bf97e4",
   955 => x"87f106ab",
   956 => x"97e4fdc0",
   957 => x"87cf02bf",
   958 => x"7087fafb",
   959 => x"c6029949",
   960 => x"a9ecc087",
   961 => x"c087f105",
   962 => x"87e9fb4b",
   963 => x"e4fb4d70",
   964 => x"58a6c887",
   965 => x"7087defb",
   966 => x"c883c14a",
   967 => x"699749a4",
   968 => x"da05ad49",
   969 => x"49a4c987",
   970 => x"c4496997",
   971 => x"ce05a966",
   972 => x"49a4ca87",
   973 => x"aa496997",
   974 => x"c187c405",
   975 => x"c087d07e",
   976 => x"c602adec",
   977 => x"adfbc087",
   978 => x"c087c405",
   979 => x"6e7ec14b",
   980 => x"87f5fe02",
   981 => x"7387fdfa",
   982 => x"268ef848",
   983 => x"264c264d",
   984 => x"004f264b",
   985 => x"1e731e00",
   986 => x"c84bd4ff",
   987 => x"d0ff4a66",
   988 => x"78c5c848",
   989 => x"c148d4ff",
   990 => x"7b1178d4",
   991 => x"f9058ac1",
   992 => x"48d0ff87",
   993 => x"4b2678c4",
   994 => x"5e0e4f26",
   995 => x"0e5d5c5b",
   996 => x"7e7186f8",
   997 => x"eec21e6e",
   998 => x"d8e549cc",
   999 => x"7086c487",
  1000 => x"e4c40298",
  1001 => x"ececc187",
  1002 => x"496e4cbf",
  1003 => x"c887d6fc",
  1004 => x"987058a6",
  1005 => x"c487c505",
  1006 => x"78c148a6",
  1007 => x"c548d0ff",
  1008 => x"48d4ff78",
  1009 => x"c478d5c1",
  1010 => x"89c14966",
  1011 => x"ecc131c6",
  1012 => x"4abf97e4",
  1013 => x"ffb07148",
  1014 => x"ff7808d4",
  1015 => x"78c448d0",
  1016 => x"97c8eec2",
  1017 => x"99d049bf",
  1018 => x"c587dd02",
  1019 => x"48d4ff78",
  1020 => x"c078d6c1",
  1021 => x"48d4ff4a",
  1022 => x"c178ffc3",
  1023 => x"aae0c082",
  1024 => x"ff87f204",
  1025 => x"78c448d0",
  1026 => x"c348d4ff",
  1027 => x"d0ff78ff",
  1028 => x"ff78c548",
  1029 => x"d3c148d4",
  1030 => x"ff78c178",
  1031 => x"78c448d0",
  1032 => x"06acb7c0",
  1033 => x"c287cbc2",
  1034 => x"4bbfd4ee",
  1035 => x"737e748c",
  1036 => x"ddc1029b",
  1037 => x"4dc0c887",
  1038 => x"abb7c08b",
  1039 => x"c887c603",
  1040 => x"c04da3c0",
  1041 => x"c8eec24b",
  1042 => x"d049bf97",
  1043 => x"87cf0299",
  1044 => x"eec21ec0",
  1045 => x"e2e749cc",
  1046 => x"7086c487",
  1047 => x"c287d84c",
  1048 => x"c21ecce1",
  1049 => x"e749ccee",
  1050 => x"4c7087d1",
  1051 => x"e1c21e75",
  1052 => x"f0fb49cc",
  1053 => x"7486c887",
  1054 => x"87c5059c",
  1055 => x"cac148c0",
  1056 => x"c21ec187",
  1057 => x"e549ccee",
  1058 => x"86c487d2",
  1059 => x"fe059b73",
  1060 => x"4c6e87e3",
  1061 => x"06acb7c0",
  1062 => x"eec287d1",
  1063 => x"78c048cc",
  1064 => x"78c080d0",
  1065 => x"eec280f4",
  1066 => x"c078bfd8",
  1067 => x"fd01acb7",
  1068 => x"d0ff87f5",
  1069 => x"ff78c548",
  1070 => x"d3c148d4",
  1071 => x"ff78c078",
  1072 => x"78c448d0",
  1073 => x"c2c048c1",
  1074 => x"f848c087",
  1075 => x"264d268e",
  1076 => x"264b264c",
  1077 => x"5b5e0e4f",
  1078 => x"fc0e5d5c",
  1079 => x"c04d7186",
  1080 => x"04ad4c4b",
  1081 => x"c087e8c0",
  1082 => x"741ec5fb",
  1083 => x"87c4029c",
  1084 => x"87c24ac0",
  1085 => x"49724ac1",
  1086 => x"c487e0eb",
  1087 => x"c17e7086",
  1088 => x"c2056e83",
  1089 => x"c14b7587",
  1090 => x"06ab7584",
  1091 => x"6e87d8ff",
  1092 => x"268efc48",
  1093 => x"264c264d",
  1094 => x"0e4f264b",
  1095 => x"0e5c5b5e",
  1096 => x"66cc4b71",
  1097 => x"4c87d802",
  1098 => x"028cf0c0",
  1099 => x"4a7487d8",
  1100 => x"d1028ac1",
  1101 => x"cd028a87",
  1102 => x"c9028a87",
  1103 => x"7387d987",
  1104 => x"87c6f949",
  1105 => x"1e7487d2",
  1106 => x"d8c149c0",
  1107 => x"1e7487ee",
  1108 => x"d8c14973",
  1109 => x"86c887e6",
  1110 => x"4b264c26",
  1111 => x"5e0e4f26",
  1112 => x"0e5d5c5b",
  1113 => x"4c7186fc",
  1114 => x"c291de49",
  1115 => x"714df8ee",
  1116 => x"026d9785",
  1117 => x"c287dcc1",
  1118 => x"49bfe8ee",
  1119 => x"fd718174",
  1120 => x"7e7087d3",
  1121 => x"c0029848",
  1122 => x"eec287f2",
  1123 => x"4a704bec",
  1124 => x"fefe49cb",
  1125 => x"4b7487ce",
  1126 => x"ecc193cc",
  1127 => x"83c483f0",
  1128 => x"7be0c7c1",
  1129 => x"c3c14974",
  1130 => x"7b7587de",
  1131 => x"97e8ecc1",
  1132 => x"c21e49bf",
  1133 => x"fd49ecee",
  1134 => x"86c487e1",
  1135 => x"c3c14974",
  1136 => x"49c087c6",
  1137 => x"87e1c4c1",
  1138 => x"48c4eec2",
  1139 => x"c04950c0",
  1140 => x"fc87cce2",
  1141 => x"264d268e",
  1142 => x"264b264c",
  1143 => x"0000004f",
  1144 => x"64616f4c",
  1145 => x"2e676e69",
  1146 => x"1e002e2e",
  1147 => x"4b711e73",
  1148 => x"e8eec249",
  1149 => x"fb7181bf",
  1150 => x"4a7087db",
  1151 => x"87c4029a",
  1152 => x"87dde649",
  1153 => x"48e8eec2",
  1154 => x"497378c0",
  1155 => x"2687fac1",
  1156 => x"1e4f264b",
  1157 => x"4b711e73",
  1158 => x"024aa3c4",
  1159 => x"c187d0c1",
  1160 => x"87dc028a",
  1161 => x"f2c0028a",
  1162 => x"c1058a87",
  1163 => x"eec287d3",
  1164 => x"c102bfe8",
  1165 => x"c14887cb",
  1166 => x"eceec288",
  1167 => x"87c1c158",
  1168 => x"bfe8eec2",
  1169 => x"c289c649",
  1170 => x"c059ecee",
  1171 => x"c003a9b7",
  1172 => x"eec287ef",
  1173 => x"78c048e8",
  1174 => x"c287e6c0",
  1175 => x"02bfe4ee",
  1176 => x"eec287df",
  1177 => x"c148bfe8",
  1178 => x"eceec280",
  1179 => x"c287d258",
  1180 => x"02bfe4ee",
  1181 => x"eec287cb",
  1182 => x"c648bfe8",
  1183 => x"eceec280",
  1184 => x"c4497358",
  1185 => x"264b2687",
  1186 => x"5b5e0e4f",
  1187 => x"f00e5d5c",
  1188 => x"59a6d086",
  1189 => x"4dcce1c2",
  1190 => x"eec24cc0",
  1191 => x"78c148e4",
  1192 => x"c048a6c4",
  1193 => x"c27e7578",
  1194 => x"48bfe8ee",
  1195 => x"c006a8c0",
  1196 => x"7e7587fa",
  1197 => x"48cce1c2",
  1198 => x"efc00298",
  1199 => x"c5fbc087",
  1200 => x"0266c81e",
  1201 => x"4dc087c4",
  1202 => x"4dc187c2",
  1203 => x"cae44975",
  1204 => x"7086c487",
  1205 => x"c484c17e",
  1206 => x"80c14866",
  1207 => x"c258a6c8",
  1208 => x"acbfe8ee",
  1209 => x"6e87c503",
  1210 => x"87d1ff05",
  1211 => x"4cc04d6e",
  1212 => x"c3029d75",
  1213 => x"fbc087e0",
  1214 => x"66c81ec5",
  1215 => x"cc87c702",
  1216 => x"78c048a6",
  1217 => x"a6cc87c5",
  1218 => x"cc78c148",
  1219 => x"cae34966",
  1220 => x"7086c487",
  1221 => x"0298487e",
  1222 => x"4987e8c2",
  1223 => x"699781cb",
  1224 => x"0299d049",
  1225 => x"c187d6c1",
  1226 => x"744aebc7",
  1227 => x"c191cc49",
  1228 => x"7281f0ec",
  1229 => x"c381c879",
  1230 => x"497451ff",
  1231 => x"eec291de",
  1232 => x"85714df8",
  1233 => x"7d97c1c2",
  1234 => x"c049a5c1",
  1235 => x"e9c251e0",
  1236 => x"02bf97dc",
  1237 => x"84c187d2",
  1238 => x"c24ba5c2",
  1239 => x"db4adce9",
  1240 => x"fff6fe49",
  1241 => x"87dbc187",
  1242 => x"c049a5cd",
  1243 => x"c284c151",
  1244 => x"4a6e4ba5",
  1245 => x"f6fe49cb",
  1246 => x"c6c187ea",
  1247 => x"dec5c187",
  1248 => x"cc49744a",
  1249 => x"f0ecc191",
  1250 => x"c2797281",
  1251 => x"bf97dce9",
  1252 => x"7487d802",
  1253 => x"c191de49",
  1254 => x"f8eec284",
  1255 => x"c283714b",
  1256 => x"dd4adce9",
  1257 => x"fbf5fe49",
  1258 => x"7487d887",
  1259 => x"c293de4b",
  1260 => x"cb83f8ee",
  1261 => x"51c049a3",
  1262 => x"6e7384c1",
  1263 => x"fe49cb4a",
  1264 => x"c487e1f5",
  1265 => x"80c14866",
  1266 => x"c758a6c8",
  1267 => x"c5c003ac",
  1268 => x"fc056e87",
  1269 => x"acc787e0",
  1270 => x"87e6c003",
  1271 => x"48e4eec2",
  1272 => x"c5c178c0",
  1273 => x"49744ade",
  1274 => x"ecc191cc",
  1275 => x"797281f0",
  1276 => x"91de4974",
  1277 => x"81f8eec2",
  1278 => x"84c151c0",
  1279 => x"ff04acc7",
  1280 => x"eec187da",
  1281 => x"50c048cc",
  1282 => x"d1c180f7",
  1283 => x"d0c140f9",
  1284 => x"80c878ec",
  1285 => x"78d3c8c1",
  1286 => x"c04966cc",
  1287 => x"f087e9f9",
  1288 => x"264d268e",
  1289 => x"264b264c",
  1290 => x"0000004f",
  1291 => x"61422080",
  1292 => x"1e006b63",
  1293 => x"4b711e73",
  1294 => x"c191cc49",
  1295 => x"c881f0ec",
  1296 => x"ecc14aa1",
  1297 => x"501248e4",
  1298 => x"c04aa1c9",
  1299 => x"1248e4fd",
  1300 => x"c181ca50",
  1301 => x"1148e8ec",
  1302 => x"e8ecc150",
  1303 => x"1e49bf97",
  1304 => x"f6f249c0",
  1305 => x"f8497387",
  1306 => x"8efc87df",
  1307 => x"4f264b26",
  1308 => x"c049c01e",
  1309 => x"2687f2f9",
  1310 => x"4a711e4f",
  1311 => x"c191cc49",
  1312 => x"c881f0ec",
  1313 => x"c4eec281",
  1314 => x"c0501148",
  1315 => x"fe49a2f0",
  1316 => x"c087f9ef",
  1317 => x"87c7d749",
  1318 => x"ff1e4f26",
  1319 => x"ffc34ad4",
  1320 => x"48d0ff7a",
  1321 => x"de78e1c0",
  1322 => x"487a717a",
  1323 => x"7028b7c8",
  1324 => x"d048717a",
  1325 => x"7a7028b7",
  1326 => x"b7d84871",
  1327 => x"ff7a7028",
  1328 => x"e0c048d0",
  1329 => x"0e4f2678",
  1330 => x"5d5c5b5e",
  1331 => x"7186f40e",
  1332 => x"91cc494d",
  1333 => x"81f0ecc1",
  1334 => x"ca4aa1c8",
  1335 => x"a6c47ea1",
  1336 => x"c0eec248",
  1337 => x"976e78bf",
  1338 => x"66c44bbf",
  1339 => x"122c734c",
  1340 => x"58a6cc48",
  1341 => x"84c19c70",
  1342 => x"699781c9",
  1343 => x"04acb749",
  1344 => x"4cc087c2",
  1345 => x"4abf976e",
  1346 => x"724966c8",
  1347 => x"c4b9ff31",
  1348 => x"48749966",
  1349 => x"4a703072",
  1350 => x"c4eec2b1",
  1351 => x"f9fd7159",
  1352 => x"c21ec787",
  1353 => x"1ebfe0ee",
  1354 => x"1ef0ecc1",
  1355 => x"97c4eec2",
  1356 => x"f4c149bf",
  1357 => x"c0497587",
  1358 => x"e887cdf5",
  1359 => x"264d268e",
  1360 => x"264b264c",
  1361 => x"1e731e4f",
  1362 => x"fd494b71",
  1363 => x"497387f9",
  1364 => x"2687f4fd",
  1365 => x"1e4f264b",
  1366 => x"4b711e73",
  1367 => x"024aa3c2",
  1368 => x"8ac187d6",
  1369 => x"87e2c005",
  1370 => x"bfe0eec2",
  1371 => x"4887db02",
  1372 => x"eec288c1",
  1373 => x"87d258e4",
  1374 => x"bfe4eec2",
  1375 => x"c287cb02",
  1376 => x"48bfe0ee",
  1377 => x"eec280c1",
  1378 => x"1ec758e4",
  1379 => x"bfe0eec2",
  1380 => x"f0ecc11e",
  1381 => x"c4eec21e",
  1382 => x"cc49bf97",
  1383 => x"c0497387",
  1384 => x"f487e5f3",
  1385 => x"264b268e",
  1386 => x"5b5e0e4f",
  1387 => x"ff0e5d5c",
  1388 => x"e4c086cc",
  1389 => x"a6cc59a6",
  1390 => x"c478c048",
  1391 => x"c478c080",
  1392 => x"66c8c180",
  1393 => x"c180c478",
  1394 => x"c180c478",
  1395 => x"e4eec278",
  1396 => x"e078c148",
  1397 => x"c4e187ea",
  1398 => x"87d9e087",
  1399 => x"fbc04c70",
  1400 => x"f3c102ac",
  1401 => x"66e0c087",
  1402 => x"87e8c105",
  1403 => x"4a66c4c1",
  1404 => x"7e6a82c4",
  1405 => x"48c0e9c1",
  1406 => x"4120496e",
  1407 => x"51104120",
  1408 => x"4866c4c1",
  1409 => x"78f3d0c1",
  1410 => x"81c7496a",
  1411 => x"c4c15174",
  1412 => x"81c84966",
  1413 => x"a6d851c1",
  1414 => x"c178c248",
  1415 => x"c94966c4",
  1416 => x"c151c081",
  1417 => x"ca4966c4",
  1418 => x"c151c081",
  1419 => x"6a1ed81e",
  1420 => x"ff81c849",
  1421 => x"c887fadf",
  1422 => x"66c8c186",
  1423 => x"01a8c048",
  1424 => x"a6d087c7",
  1425 => x"cf78c148",
  1426 => x"66c8c187",
  1427 => x"d888c148",
  1428 => x"87c458a6",
  1429 => x"87c5dfff",
  1430 => x"cd029c74",
  1431 => x"66d087da",
  1432 => x"66ccc148",
  1433 => x"cfcd03a8",
  1434 => x"48a6c887",
  1435 => x"ff7e78c0",
  1436 => x"7087c2de",
  1437 => x"acd0c14c",
  1438 => x"87e7c205",
  1439 => x"6e48a6c4",
  1440 => x"87d8e078",
  1441 => x"cc487e70",
  1442 => x"c506a866",
  1443 => x"48a6cc87",
  1444 => x"ddff786e",
  1445 => x"4c7087df",
  1446 => x"05acecc0",
  1447 => x"d087eec1",
  1448 => x"91cc4966",
  1449 => x"8166c4c1",
  1450 => x"6a4aa1c4",
  1451 => x"4aa1c84d",
  1452 => x"d1c1526e",
  1453 => x"dcff79f9",
  1454 => x"4c7087fb",
  1455 => x"87d9029c",
  1456 => x"02acfbc0",
  1457 => x"557487d3",
  1458 => x"87e9dcff",
  1459 => x"029c4c70",
  1460 => x"fbc087c7",
  1461 => x"edff05ac",
  1462 => x"55e0c087",
  1463 => x"c055c1c2",
  1464 => x"e0c07d97",
  1465 => x"66c44866",
  1466 => x"87db05a8",
  1467 => x"d44866d0",
  1468 => x"ca04a866",
  1469 => x"4866d087",
  1470 => x"a6d480c1",
  1471 => x"d487c858",
  1472 => x"88c14866",
  1473 => x"ff58a6d8",
  1474 => x"7087eadb",
  1475 => x"acd0c14c",
  1476 => x"dc87c905",
  1477 => x"80c14866",
  1478 => x"58a6e0c0",
  1479 => x"02acd0c1",
  1480 => x"6e87d9fd",
  1481 => x"66e0c048",
  1482 => x"ebc905a8",
  1483 => x"a6e4c087",
  1484 => x"7478c048",
  1485 => x"88fbc048",
  1486 => x"7058a6c8",
  1487 => x"ddc90298",
  1488 => x"88cb4887",
  1489 => x"7058a6c8",
  1490 => x"cfc10298",
  1491 => x"88c94887",
  1492 => x"7058a6c8",
  1493 => x"ffc30298",
  1494 => x"88c44887",
  1495 => x"7058a6c8",
  1496 => x"87cf0298",
  1497 => x"c888c148",
  1498 => x"987058a6",
  1499 => x"87e8c302",
  1500 => x"c887dcc8",
  1501 => x"f0c048a6",
  1502 => x"f8d9ff78",
  1503 => x"c04c7087",
  1504 => x"c002acec",
  1505 => x"a6cc87c3",
  1506 => x"acecc05c",
  1507 => x"ff87cd02",
  1508 => x"7087e2d9",
  1509 => x"acecc04c",
  1510 => x"87f3ff05",
  1511 => x"02acecc0",
  1512 => x"ff87c4c0",
  1513 => x"c087ced9",
  1514 => x"d81eca1e",
  1515 => x"91cc4966",
  1516 => x"4866ccc1",
  1517 => x"a6cc8071",
  1518 => x"4866c858",
  1519 => x"a6d080c4",
  1520 => x"bf66cc58",
  1521 => x"e8d9ff49",
  1522 => x"de1ec187",
  1523 => x"bf66d41e",
  1524 => x"dcd9ff49",
  1525 => x"7086d087",
  1526 => x"08c04849",
  1527 => x"a6ecc088",
  1528 => x"06a8c058",
  1529 => x"c087eec0",
  1530 => x"dd4866e8",
  1531 => x"e4c003a8",
  1532 => x"bf66c487",
  1533 => x"66e8c049",
  1534 => x"51e0c081",
  1535 => x"4966e8c0",
  1536 => x"66c481c1",
  1537 => x"c1c281bf",
  1538 => x"66e8c051",
  1539 => x"c481c249",
  1540 => x"c081bf66",
  1541 => x"c1486e51",
  1542 => x"6e78f3d0",
  1543 => x"d881c849",
  1544 => x"496e5166",
  1545 => x"66dc81c9",
  1546 => x"ca496e51",
  1547 => x"5166c881",
  1548 => x"c14866d8",
  1549 => x"58a6dc80",
  1550 => x"d44866d0",
  1551 => x"c004a866",
  1552 => x"66d087cb",
  1553 => x"d480c148",
  1554 => x"d1c558a6",
  1555 => x"4866d487",
  1556 => x"a6d888c1",
  1557 => x"87c6c558",
  1558 => x"87c0d9ff",
  1559 => x"58a6ecc0",
  1560 => x"87f8d8ff",
  1561 => x"58a6f0c0",
  1562 => x"05a8ecc0",
  1563 => x"a687c9c0",
  1564 => x"66e8c048",
  1565 => x"87c4c078",
  1566 => x"87f9d5ff",
  1567 => x"cc4966d0",
  1568 => x"66c4c191",
  1569 => x"c8807148",
  1570 => x"66c458a6",
  1571 => x"c482c84a",
  1572 => x"81ca4966",
  1573 => x"5166e8c0",
  1574 => x"4966ecc0",
  1575 => x"e8c081c1",
  1576 => x"48c18966",
  1577 => x"49703071",
  1578 => x"977189c1",
  1579 => x"c0eec27a",
  1580 => x"e8c049bf",
  1581 => x"6a972966",
  1582 => x"9871484a",
  1583 => x"58a6f4c0",
  1584 => x"c44866c4",
  1585 => x"58a6cc80",
  1586 => x"4dbf66c8",
  1587 => x"4866e0c0",
  1588 => x"c002a86e",
  1589 => x"7ec087c5",
  1590 => x"c187c2c0",
  1591 => x"c01e6e7e",
  1592 => x"49751ee0",
  1593 => x"87c9d5ff",
  1594 => x"4c7086c8",
  1595 => x"06acb7c0",
  1596 => x"7487d4c1",
  1597 => x"bf66c885",
  1598 => x"81e0c049",
  1599 => x"c14b8975",
  1600 => x"714acce9",
  1601 => x"87dce0fe",
  1602 => x"7e7585c2",
  1603 => x"4866e4c0",
  1604 => x"e8c080c1",
  1605 => x"f0c058a6",
  1606 => x"81c14966",
  1607 => x"c002a970",
  1608 => x"4dc087c5",
  1609 => x"c187c2c0",
  1610 => x"cc1e754d",
  1611 => x"c049bf66",
  1612 => x"66c481e0",
  1613 => x"c81e7189",
  1614 => x"d3ff4966",
  1615 => x"86c887f3",
  1616 => x"01a8b7c0",
  1617 => x"c087c5ff",
  1618 => x"c00266e4",
  1619 => x"66c487d3",
  1620 => x"c081c949",
  1621 => x"c45166e4",
  1622 => x"d3c14866",
  1623 => x"cec078c7",
  1624 => x"4966c487",
  1625 => x"51c281c9",
  1626 => x"c14866c4",
  1627 => x"d078c5d5",
  1628 => x"66d44866",
  1629 => x"cbc004a8",
  1630 => x"4866d087",
  1631 => x"a6d480c1",
  1632 => x"87dac058",
  1633 => x"c14866d4",
  1634 => x"58a6d888",
  1635 => x"ff87cfc0",
  1636 => x"7087cad2",
  1637 => x"87c6c04c",
  1638 => x"87c1d2ff",
  1639 => x"66dc4c70",
  1640 => x"c080c148",
  1641 => x"7458a6e0",
  1642 => x"cbc0029c",
  1643 => x"4866d087",
  1644 => x"a866ccc1",
  1645 => x"87f1f204",
  1646 => x"c74866d0",
  1647 => x"e1c003a8",
  1648 => x"4c66d087",
  1649 => x"48e4eec2",
  1650 => x"497478c0",
  1651 => x"c4c191cc",
  1652 => x"a1c48166",
  1653 => x"c04a6a4a",
  1654 => x"84c17952",
  1655 => x"ff04acc7",
  1656 => x"e0c087e2",
  1657 => x"e2c00266",
  1658 => x"66c4c187",
  1659 => x"81d4c149",
  1660 => x"4a66c4c1",
  1661 => x"c082dcc1",
  1662 => x"f9d1c152",
  1663 => x"66c4c179",
  1664 => x"81d8c149",
  1665 => x"79d0e9c1",
  1666 => x"c187d6c0",
  1667 => x"c14966c4",
  1668 => x"c4c181d4",
  1669 => x"d8c14a66",
  1670 => x"d8e9c182",
  1671 => x"f0d1c17a",
  1672 => x"d7d5c179",
  1673 => x"66c4c14a",
  1674 => x"81e0c149",
  1675 => x"cfff7972",
  1676 => x"66cc87e2",
  1677 => x"8eccff48",
  1678 => x"4c264d26",
  1679 => x"4f264b26",
  1680 => x"64616f4c",
  1681 => x"202e2a20",
  1682 => x"00000000",
  1683 => x"0000203a",
  1684 => x"61422080",
  1685 => x"00006b63",
  1686 => x"78452080",
  1687 => x"1e007469",
  1688 => x"eec21ec7",
  1689 => x"c11ebfe0",
  1690 => x"c21ef0ec",
  1691 => x"bf97c4ee",
  1692 => x"87f5ec49",
  1693 => x"49f0ecc1",
  1694 => x"87dae1c0",
  1695 => x"4f268ef4",
  1696 => x"c81e731e",
  1697 => x"eec287c3",
  1698 => x"50c048ec",
  1699 => x"48c8eec1",
  1700 => x"78d0ecc1",
  1701 => x"49a0e8fe",
  1702 => x"87fae0c0",
  1703 => x"e7df49c7",
  1704 => x"c049c187",
  1705 => x"ff87c2e1",
  1706 => x"ffc348d4",
  1707 => x"dbe3fe78",
  1708 => x"02987087",
  1709 => x"edfe87cd",
  1710 => x"987087d7",
  1711 => x"c187c402",
  1712 => x"c087c24a",
  1713 => x"029a724a",
  1714 => x"ecc187c8",
  1715 => x"d7fe49dc",
  1716 => x"eec287d5",
  1717 => x"78c048e0",
  1718 => x"48c4eec2",
  1719 => x"fd4950c0",
  1720 => x"f4c087fd",
  1721 => x"4b7087da",
  1722 => x"87cb029b",
  1723 => x"5bcceec1",
  1724 => x"d3de49c7",
  1725 => x"c087c587",
  1726 => x"87eddf49",
  1727 => x"c087c4c3",
  1728 => x"c087cee1",
  1729 => x"ff87e2ee",
  1730 => x"4b2687f5",
  1731 => x"00004f26",
  1732 => x"746f6f42",
  1733 => x"2e676e69",
  1734 => x"00002e2e",
  1735 => x"4f204453",
  1736 => x"0000004b",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"00000001",
  1740 => x"0000115e",
  1741 => x"00002bb8",
  1742 => x"00000000",
  1743 => x"0000115e",
  1744 => x"00002bd6",
  1745 => x"00000000",
  1746 => x"0000115e",
  1747 => x"00002bf4",
  1748 => x"00000000",
  1749 => x"0000115e",
  1750 => x"00002c12",
  1751 => x"00000000",
  1752 => x"0000115e",
  1753 => x"00002c30",
  1754 => x"00000000",
  1755 => x"0000115e",
  1756 => x"00002c4e",
  1757 => x"00000000",
  1758 => x"0000115e",
  1759 => x"00002c6c",
  1760 => x"00000000",
  1761 => x"00001479",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00001213",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"db86fc1e",
  1768 => x"fc7e7087",
  1769 => x"1e4f268e",
  1770 => x"c048f0fe",
  1771 => x"7909cd78",
  1772 => x"1e4f2609",
  1773 => x"49dceec1",
  1774 => x"4f2687ed",
  1775 => x"bff0fe1e",
  1776 => x"1e4f2648",
  1777 => x"c148f0fe",
  1778 => x"1e4f2678",
  1779 => x"c048f0fe",
  1780 => x"1e4f2678",
  1781 => x"52c04a71",
  1782 => x"0e4f2651",
  1783 => x"5d5c5b5e",
  1784 => x"7186f40e",
  1785 => x"7e6d974d",
  1786 => x"974ca5c1",
  1787 => x"a6c8486c",
  1788 => x"c4486e58",
  1789 => x"c505a866",
  1790 => x"c048ff87",
  1791 => x"caff87e6",
  1792 => x"49a5c287",
  1793 => x"714b6c97",
  1794 => x"6b974ba3",
  1795 => x"7e6c974b",
  1796 => x"80c1486e",
  1797 => x"c758a6c8",
  1798 => x"58a6cc98",
  1799 => x"fe7c9770",
  1800 => x"487387e1",
  1801 => x"4d268ef4",
  1802 => x"4b264c26",
  1803 => x"5e0e4f26",
  1804 => x"f40e5c5b",
  1805 => x"d84c7186",
  1806 => x"ffc34a66",
  1807 => x"4ba4c29a",
  1808 => x"73496c97",
  1809 => x"517249a1",
  1810 => x"6e7e6c97",
  1811 => x"c880c148",
  1812 => x"98c758a6",
  1813 => x"7058a6cc",
  1814 => x"268ef454",
  1815 => x"264b264c",
  1816 => x"86fc1e4f",
  1817 => x"e087e4fd",
  1818 => x"c0494abf",
  1819 => x"0299c0e0",
  1820 => x"1e7287cb",
  1821 => x"49ccf2c2",
  1822 => x"c487f3fe",
  1823 => x"87fcfc86",
  1824 => x"fefc7e70",
  1825 => x"268efc87",
  1826 => x"f2c21e4f",
  1827 => x"c2fd49cc",
  1828 => x"e1f1c187",
  1829 => x"87cffc49",
  1830 => x"2687f1c2",
  1831 => x"1e731e4f",
  1832 => x"49ccf2c2",
  1833 => x"7087f4fc",
  1834 => x"aab7c04a",
  1835 => x"87ccc204",
  1836 => x"05aaf0c3",
  1837 => x"f5c187c9",
  1838 => x"78c148c4",
  1839 => x"c387edc1",
  1840 => x"c905aae0",
  1841 => x"c8f5c187",
  1842 => x"c178c148",
  1843 => x"f5c187de",
  1844 => x"c602bfc8",
  1845 => x"a2c0c287",
  1846 => x"7287c24b",
  1847 => x"c4f5c14b",
  1848 => x"e0c002bf",
  1849 => x"c4497387",
  1850 => x"c19129b7",
  1851 => x"7381e0f6",
  1852 => x"c29acf4a",
  1853 => x"7248c192",
  1854 => x"ff4a7030",
  1855 => x"694872ba",
  1856 => x"db797098",
  1857 => x"c4497387",
  1858 => x"c19129b7",
  1859 => x"7381e0f6",
  1860 => x"c29acf4a",
  1861 => x"7248c392",
  1862 => x"484a7030",
  1863 => x"7970b069",
  1864 => x"48c8f5c1",
  1865 => x"f5c178c0",
  1866 => x"78c048c4",
  1867 => x"49ccf2c2",
  1868 => x"7087e8fa",
  1869 => x"aab7c04a",
  1870 => x"87f4fd03",
  1871 => x"4b2648c0",
  1872 => x"00004f26",
  1873 => x"00000000",
  1874 => x"00000000",
  1875 => x"724ac01e",
  1876 => x"c191c449",
  1877 => x"c081e0f6",
  1878 => x"d082c179",
  1879 => x"ee04aab7",
  1880 => x"0e4f2687",
  1881 => x"5d5c5b5e",
  1882 => x"f94d710e",
  1883 => x"4a7587dd",
  1884 => x"922ab7c4",
  1885 => x"82e0f6c1",
  1886 => x"9ccf4c75",
  1887 => x"496a94c2",
  1888 => x"c32b744b",
  1889 => x"7448c29b",
  1890 => x"ff4c7030",
  1891 => x"714874bc",
  1892 => x"f87a7098",
  1893 => x"487387ed",
  1894 => x"4c264d26",
  1895 => x"4f264b26",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"48d0ff1e",
  1913 => x"7178e1c8",
  1914 => x"08d4ff48",
  1915 => x"1e4f2678",
  1916 => x"c848d0ff",
  1917 => x"487178e1",
  1918 => x"7808d4ff",
  1919 => x"ff4866c4",
  1920 => x"267808d4",
  1921 => x"4a711e4f",
  1922 => x"1e4966c4",
  1923 => x"deff4972",
  1924 => x"48d0ff87",
  1925 => x"fc78e0c0",
  1926 => x"1e4f268e",
  1927 => x"4b711e73",
  1928 => x"1e4966c8",
  1929 => x"e0c14a73",
  1930 => x"d8ff49a2",
  1931 => x"268efc87",
  1932 => x"1e4f264b",
  1933 => x"c848d0ff",
  1934 => x"487178c9",
  1935 => x"7808d4ff",
  1936 => x"711e4f26",
  1937 => x"87eb494a",
  1938 => x"c848d0ff",
  1939 => x"1e4f2678",
  1940 => x"4b711e73",
  1941 => x"bfe4f2c2",
  1942 => x"c287c302",
  1943 => x"d0ff87eb",
  1944 => x"78c9c848",
  1945 => x"e0c04873",
  1946 => x"08d4ffb0",
  1947 => x"d8f2c278",
  1948 => x"c878c048",
  1949 => x"87c50266",
  1950 => x"c249ffc3",
  1951 => x"c249c087",
  1952 => x"cc59e0f2",
  1953 => x"87c60266",
  1954 => x"4ad5d5c5",
  1955 => x"ffcf87c4",
  1956 => x"f2c24aff",
  1957 => x"f2c25ae4",
  1958 => x"78c148e4",
  1959 => x"4f264b26",
  1960 => x"5c5b5e0e",
  1961 => x"4d710e5d",
  1962 => x"bfe0f2c2",
  1963 => x"029d754b",
  1964 => x"c84987cb",
  1965 => x"c8f9c191",
  1966 => x"c482714a",
  1967 => x"c8fdc187",
  1968 => x"124cc04a",
  1969 => x"c2997349",
  1970 => x"48bfdcf2",
  1971 => x"d4ffb871",
  1972 => x"b7c17808",
  1973 => x"b7c8842b",
  1974 => x"87e704ac",
  1975 => x"bfd8f2c2",
  1976 => x"c280c848",
  1977 => x"2658dcf2",
  1978 => x"264c264d",
  1979 => x"1e4f264b",
  1980 => x"4b711e73",
  1981 => x"029a4a13",
  1982 => x"497287cb",
  1983 => x"1387e1fe",
  1984 => x"f5059a4a",
  1985 => x"264b2687",
  1986 => x"f2c21e4f",
  1987 => x"c249bfd8",
  1988 => x"c148d8f2",
  1989 => x"c0c478a1",
  1990 => x"db03a9b7",
  1991 => x"48d4ff87",
  1992 => x"bfdcf2c2",
  1993 => x"d8f2c278",
  1994 => x"f2c249bf",
  1995 => x"a1c148d8",
  1996 => x"b7c0c478",
  1997 => x"87e504a9",
  1998 => x"c848d0ff",
  1999 => x"e4f2c278",
  2000 => x"2678c048",
  2001 => x"0000004f",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"5f000000",
  2005 => x"0000005f",
  2006 => x"00030300",
  2007 => x"00000303",
  2008 => x"147f7f14",
  2009 => x"00147f7f",
  2010 => x"6b2e2400",
  2011 => x"00123a6b",
  2012 => x"18366a4c",
  2013 => x"0032566c",
  2014 => x"594f7e30",
  2015 => x"40683a77",
  2016 => x"07040000",
  2017 => x"00000003",
  2018 => x"3e1c0000",
  2019 => x"00004163",
  2020 => x"63410000",
  2021 => x"00001c3e",
  2022 => x"1c3e2a08",
  2023 => x"082a3e1c",
  2024 => x"3e080800",
  2025 => x"0008083e",
  2026 => x"e0800000",
  2027 => x"00000060",
  2028 => x"08080800",
  2029 => x"00080808",
  2030 => x"60000000",
  2031 => x"00000060",
  2032 => x"18306040",
  2033 => x"0103060c",
  2034 => x"597f3e00",
  2035 => x"003e7f4d",
  2036 => x"7f060400",
  2037 => x"0000007f",
  2038 => x"71634200",
  2039 => x"00464f59",
  2040 => x"49632200",
  2041 => x"00367f49",
  2042 => x"13161c18",
  2043 => x"00107f7f",
  2044 => x"45672700",
  2045 => x"00397d45",
  2046 => x"4b7e3c00",
  2047 => x"00307949",
  2048 => x"71010100",
  2049 => x"00070f79",
  2050 => x"497f3600",
  2051 => x"00367f49",
  2052 => x"494f0600",
  2053 => x"001e3f69",
  2054 => x"66000000",
  2055 => x"00000066",
  2056 => x"e6800000",
  2057 => x"00000066",
  2058 => x"14080800",
  2059 => x"00222214",
  2060 => x"14141400",
  2061 => x"00141414",
  2062 => x"14222200",
  2063 => x"00080814",
  2064 => x"51030200",
  2065 => x"00060f59",
  2066 => x"5d417f3e",
  2067 => x"001e1f55",
  2068 => x"097f7e00",
  2069 => x"007e7f09",
  2070 => x"497f7f00",
  2071 => x"00367f49",
  2072 => x"633e1c00",
  2073 => x"00414141",
  2074 => x"417f7f00",
  2075 => x"001c3e63",
  2076 => x"497f7f00",
  2077 => x"00414149",
  2078 => x"097f7f00",
  2079 => x"00010109",
  2080 => x"417f3e00",
  2081 => x"007a7b49",
  2082 => x"087f7f00",
  2083 => x"007f7f08",
  2084 => x"7f410000",
  2085 => x"0000417f",
  2086 => x"40602000",
  2087 => x"003f7f40",
  2088 => x"1c087f7f",
  2089 => x"00416336",
  2090 => x"407f7f00",
  2091 => x"00404040",
  2092 => x"0c067f7f",
  2093 => x"007f7f06",
  2094 => x"0c067f7f",
  2095 => x"007f7f18",
  2096 => x"417f3e00",
  2097 => x"003e7f41",
  2098 => x"097f7f00",
  2099 => x"00060f09",
  2100 => x"61417f3e",
  2101 => x"00407e7f",
  2102 => x"097f7f00",
  2103 => x"00667f19",
  2104 => x"4d6f2600",
  2105 => x"00327b59",
  2106 => x"7f010100",
  2107 => x"0001017f",
  2108 => x"407f3f00",
  2109 => x"003f7f40",
  2110 => x"703f0f00",
  2111 => x"000f3f70",
  2112 => x"18307f7f",
  2113 => x"007f7f30",
  2114 => x"1c366341",
  2115 => x"4163361c",
  2116 => x"7c060301",
  2117 => x"0103067c",
  2118 => x"4d597161",
  2119 => x"00414347",
  2120 => x"7f7f0000",
  2121 => x"00004141",
  2122 => x"0c060301",
  2123 => x"40603018",
  2124 => x"41410000",
  2125 => x"00007f7f",
  2126 => x"03060c08",
  2127 => x"00080c06",
  2128 => x"80808080",
  2129 => x"00808080",
  2130 => x"03000000",
  2131 => x"00000407",
  2132 => x"54742000",
  2133 => x"00787c54",
  2134 => x"447f7f00",
  2135 => x"00387c44",
  2136 => x"447c3800",
  2137 => x"00004444",
  2138 => x"447c3800",
  2139 => x"007f7f44",
  2140 => x"547c3800",
  2141 => x"00185c54",
  2142 => x"7f7e0400",
  2143 => x"00000505",
  2144 => x"a4bc1800",
  2145 => x"007cfca4",
  2146 => x"047f7f00",
  2147 => x"00787c04",
  2148 => x"3d000000",
  2149 => x"0000407d",
  2150 => x"80808000",
  2151 => x"00007dfd",
  2152 => x"107f7f00",
  2153 => x"00446c38",
  2154 => x"3f000000",
  2155 => x"0000407f",
  2156 => x"180c7c7c",
  2157 => x"00787c0c",
  2158 => x"047c7c00",
  2159 => x"00787c04",
  2160 => x"447c3800",
  2161 => x"00387c44",
  2162 => x"24fcfc00",
  2163 => x"00183c24",
  2164 => x"243c1800",
  2165 => x"00fcfc24",
  2166 => x"047c7c00",
  2167 => x"00080c04",
  2168 => x"545c4800",
  2169 => x"00207454",
  2170 => x"7f3f0400",
  2171 => x"00004444",
  2172 => x"407c3c00",
  2173 => x"007c7c40",
  2174 => x"603c1c00",
  2175 => x"001c3c60",
  2176 => x"30607c3c",
  2177 => x"003c7c60",
  2178 => x"10386c44",
  2179 => x"00446c38",
  2180 => x"e0bc1c00",
  2181 => x"001c3c60",
  2182 => x"74644400",
  2183 => x"00444c5c",
  2184 => x"3e080800",
  2185 => x"00414177",
  2186 => x"7f000000",
  2187 => x"0000007f",
  2188 => x"77414100",
  2189 => x"0008083e",
  2190 => x"03010102",
  2191 => x"00010202",
  2192 => x"7f7f7f7f",
  2193 => x"007f7f7f",
  2194 => x"1c1c0808",
  2195 => x"7f7f3e3e",
  2196 => x"3e3e7f7f",
  2197 => x"08081c1c",
  2198 => x"7c181000",
  2199 => x"0010187c",
  2200 => x"7c301000",
  2201 => x"0010307c",
  2202 => x"60603010",
  2203 => x"00061e78",
  2204 => x"183c6642",
  2205 => x"0042663c",
  2206 => x"c26a3878",
  2207 => x"00386cc6",
  2208 => x"60000060",
  2209 => x"00600000",
  2210 => x"5c5b5e0e",
  2211 => x"86fc0e5d",
  2212 => x"f2c27e71",
  2213 => x"c04cbfec",
  2214 => x"c41ec04b",
  2215 => x"c402ab66",
  2216 => x"c24dc087",
  2217 => x"754dc187",
  2218 => x"ee49731e",
  2219 => x"86c887e1",
  2220 => x"ef49e0c0",
  2221 => x"a4c487ea",
  2222 => x"f0496a4a",
  2223 => x"c8f187f1",
  2224 => x"c184cc87",
  2225 => x"abb7c883",
  2226 => x"87cdff04",
  2227 => x"4d268efc",
  2228 => x"4b264c26",
  2229 => x"711e4f26",
  2230 => x"f0f2c24a",
  2231 => x"f0f2c25a",
  2232 => x"4978c748",
  2233 => x"2687e1fe",
  2234 => x"1e731e4f",
  2235 => x"b7c04a71",
  2236 => x"87d303aa",
  2237 => x"bfccd8c2",
  2238 => x"c187c405",
  2239 => x"c087c24b",
  2240 => x"d0d8c24b",
  2241 => x"c287c45b",
  2242 => x"fc5ad0d8",
  2243 => x"ccd8c248",
  2244 => x"c14a78bf",
  2245 => x"a2c0c19a",
  2246 => x"87e6ec49",
  2247 => x"4f264b26",
  2248 => x"c44a711e",
  2249 => x"49721e66",
  2250 => x"fc87f0eb",
  2251 => x"1e4f268e",
  2252 => x"c348d4ff",
  2253 => x"d0ff78ff",
  2254 => x"78e1c048",
  2255 => x"c148d4ff",
  2256 => x"c4487178",
  2257 => x"08d4ff30",
  2258 => x"48d0ff78",
  2259 => x"2678e0c0",
  2260 => x"5b5e0e4f",
  2261 => x"f00e5d5c",
  2262 => x"48a6c886",
  2263 => x"ec4d78c0",
  2264 => x"80fc7ebf",
  2265 => x"bfecf2c2",
  2266 => x"4cbfe878",
  2267 => x"bfccd8c2",
  2268 => x"87e9e449",
  2269 => x"ca49eecb",
  2270 => x"4b7087d6",
  2271 => x"e2e749c7",
  2272 => x"05987087",
  2273 => x"496e87c8",
  2274 => x"c10299c1",
  2275 => x"4dc187c1",
  2276 => x"c27ebfec",
  2277 => x"49bfccd8",
  2278 => x"7387c2e4",
  2279 => x"87fcc949",
  2280 => x"d7029870",
  2281 => x"c4d8c287",
  2282 => x"b9c149bf",
  2283 => x"59c8d8c2",
  2284 => x"87fbfd71",
  2285 => x"c949eecb",
  2286 => x"4b7087d6",
  2287 => x"e2e649c7",
  2288 => x"05987087",
  2289 => x"6e87c7ff",
  2290 => x"0599c149",
  2291 => x"7587fffe",
  2292 => x"e3c0029d",
  2293 => x"ccd8c287",
  2294 => x"bac14abf",
  2295 => x"5ad0d8c2",
  2296 => x"0a7a0afc",
  2297 => x"c0c19ac1",
  2298 => x"d5e949a2",
  2299 => x"49dac187",
  2300 => x"c887f0e5",
  2301 => x"78c148a6",
  2302 => x"bfccd8c2",
  2303 => x"87e9c005",
  2304 => x"ffc34974",
  2305 => x"c01e7199",
  2306 => x"87d4fc49",
  2307 => x"b7c84974",
  2308 => x"c11e7129",
  2309 => x"87c8fc49",
  2310 => x"fdc386c8",
  2311 => x"87c3e549",
  2312 => x"e449fac3",
  2313 => x"d1c787fd",
  2314 => x"c3497487",
  2315 => x"b7c899ff",
  2316 => x"74b4712c",
  2317 => x"87df029c",
  2318 => x"bfc8d8c2",
  2319 => x"87dcc749",
  2320 => x"c0059870",
  2321 => x"4cc087c4",
  2322 => x"e0c287d3",
  2323 => x"87c0c749",
  2324 => x"58ccd8c2",
  2325 => x"c287c6c0",
  2326 => x"c048c8d8",
  2327 => x"c8497478",
  2328 => x"87ce0599",
  2329 => x"e349f5c3",
  2330 => x"497087f9",
  2331 => x"c00299c2",
  2332 => x"f2c287e9",
  2333 => x"c002bff0",
  2334 => x"c14887c9",
  2335 => x"f4f2c288",
  2336 => x"c487d358",
  2337 => x"e0c14866",
  2338 => x"6e7e7080",
  2339 => x"c5c002bf",
  2340 => x"49ff4b87",
  2341 => x"a6c80f73",
  2342 => x"7478c148",
  2343 => x"0599c449",
  2344 => x"c387cec0",
  2345 => x"fae249f2",
  2346 => x"c2497087",
  2347 => x"f0c00299",
  2348 => x"f0f2c287",
  2349 => x"c7487ebf",
  2350 => x"c003a8b7",
  2351 => x"486e87cb",
  2352 => x"f2c280c1",
  2353 => x"d3c058f4",
  2354 => x"4866c487",
  2355 => x"7080e0c1",
  2356 => x"02bf6e7e",
  2357 => x"4b87c5c0",
  2358 => x"0f7349fe",
  2359 => x"c148a6c8",
  2360 => x"49fdc378",
  2361 => x"7087fce1",
  2362 => x"0299c249",
  2363 => x"c287e9c0",
  2364 => x"02bff0f2",
  2365 => x"c287c9c0",
  2366 => x"c048f0f2",
  2367 => x"87d3c078",
  2368 => x"c14866c4",
  2369 => x"7e7080e0",
  2370 => x"c002bf6e",
  2371 => x"fd4b87c5",
  2372 => x"c80f7349",
  2373 => x"78c148a6",
  2374 => x"e149fac3",
  2375 => x"497087c5",
  2376 => x"c00299c2",
  2377 => x"f2c287ea",
  2378 => x"c748bff0",
  2379 => x"c003a8b7",
  2380 => x"f2c287c9",
  2381 => x"78c748f0",
  2382 => x"c487d0c0",
  2383 => x"e0c14a66",
  2384 => x"c0026a82",
  2385 => x"fc4b87c5",
  2386 => x"c80f7349",
  2387 => x"78c148a6",
  2388 => x"f2c24dc0",
  2389 => x"50c048e8",
  2390 => x"c249eecb",
  2391 => x"4b7087f2",
  2392 => x"97e8f2c2",
  2393 => x"ddc105bf",
  2394 => x"c3497487",
  2395 => x"c00599f0",
  2396 => x"dac187cd",
  2397 => x"eadfff49",
  2398 => x"02987087",
  2399 => x"c187c7c1",
  2400 => x"4cbfe84d",
  2401 => x"99ffc349",
  2402 => x"712cb7c8",
  2403 => x"ccd8c2b4",
  2404 => x"dcff49bf",
  2405 => x"497387c7",
  2406 => x"7087c1c2",
  2407 => x"c6c00298",
  2408 => x"e8f2c287",
  2409 => x"c250c148",
  2410 => x"bf97e8f2",
  2411 => x"87d6c005",
  2412 => x"f0c34974",
  2413 => x"c6ff0599",
  2414 => x"49dac187",
  2415 => x"87e3deff",
  2416 => x"fe059870",
  2417 => x"9d7587f9",
  2418 => x"87e0c002",
  2419 => x"c248a6cc",
  2420 => x"78bff0f2",
  2421 => x"cc4966cc",
  2422 => x"4866c491",
  2423 => x"7e708071",
  2424 => x"c002bf6e",
  2425 => x"cc4b87c6",
  2426 => x"0f734966",
  2427 => x"c00266c8",
  2428 => x"f2c287c8",
  2429 => x"f249bff0",
  2430 => x"8ef087ce",
  2431 => x"4c264d26",
  2432 => x"4f264b26",
  2433 => x"00000000",
  2434 => x"00000000",
  2435 => x"00000000",
  2436 => x"ff4a711e",
  2437 => x"7249bfc8",
  2438 => x"4f2648a1",
  2439 => x"bfc8ff1e",
  2440 => x"c0c0fe89",
  2441 => x"a9c0c0c0",
  2442 => x"c087c401",
  2443 => x"c187c24a",
  2444 => x"2648724a",
  2445 => x"5b5e0e4f",
  2446 => x"710e5d5c",
  2447 => x"4cd4ff4b",
  2448 => x"c04866d0",
  2449 => x"ff49d678",
  2450 => x"c387d5de",
  2451 => x"496c7cff",
  2452 => x"7199ffc3",
  2453 => x"f0c3494d",
  2454 => x"a9e0c199",
  2455 => x"c387cb05",
  2456 => x"486c7cff",
  2457 => x"66d098c3",
  2458 => x"ffc37808",
  2459 => x"494a6c7c",
  2460 => x"ffc331c8",
  2461 => x"714a6c7c",
  2462 => x"c84972b2",
  2463 => x"7cffc331",
  2464 => x"b2714a6c",
  2465 => x"31c84972",
  2466 => x"6c7cffc3",
  2467 => x"ffb2714a",
  2468 => x"e0c048d0",
  2469 => x"029b7378",
  2470 => x"7b7287c2",
  2471 => x"4d264875",
  2472 => x"4b264c26",
  2473 => x"261e4f26",
  2474 => x"5b5e0e4f",
  2475 => x"86f80e5c",
  2476 => x"a6c81e76",
  2477 => x"87fdfd49",
  2478 => x"4b7086c4",
  2479 => x"a8c2486e",
  2480 => x"87f0c203",
  2481 => x"f0c34a73",
  2482 => x"aad0c19a",
  2483 => x"c187c702",
  2484 => x"c205aae0",
  2485 => x"497387de",
  2486 => x"c30299c8",
  2487 => x"87c6ff87",
  2488 => x"9cc34c73",
  2489 => x"c105acc2",
  2490 => x"66c487c2",
  2491 => x"7131c949",
  2492 => x"4a66c41e",
  2493 => x"f2c292d4",
  2494 => x"817249f4",
  2495 => x"87d9cffe",
  2496 => x"dbff49d8",
  2497 => x"c0c887da",
  2498 => x"cce1c21e",
  2499 => x"c6e9fd49",
  2500 => x"48d0ff87",
  2501 => x"c278e0c0",
  2502 => x"cc1ecce1",
  2503 => x"92d44a66",
  2504 => x"49f4f2c2",
  2505 => x"cdfe8172",
  2506 => x"86cc87e0",
  2507 => x"c105acc1",
  2508 => x"66c487c2",
  2509 => x"7131c949",
  2510 => x"4a66c41e",
  2511 => x"f2c292d4",
  2512 => x"817249f4",
  2513 => x"87d1cefe",
  2514 => x"1ecce1c2",
  2515 => x"d44a66c8",
  2516 => x"f4f2c292",
  2517 => x"fe817249",
  2518 => x"d787e0cb",
  2519 => x"ffd9ff49",
  2520 => x"1ec0c887",
  2521 => x"49cce1c2",
  2522 => x"87c8e7fd",
  2523 => x"d0ff86cc",
  2524 => x"78e0c048",
  2525 => x"4c268ef8",
  2526 => x"4f264b26",
  2527 => x"5c5b5e0e",
  2528 => x"86fc0e5d",
  2529 => x"d4ff4d71",
  2530 => x"7e66d44c",
  2531 => x"a8b7c348",
  2532 => x"87e2c101",
  2533 => x"66c41e75",
  2534 => x"c293d44b",
  2535 => x"7383f4f2",
  2536 => x"d0c5fe49",
  2537 => x"49a3c887",
  2538 => x"d0ff4969",
  2539 => x"78e1c848",
  2540 => x"48717cdd",
  2541 => x"7098ffc3",
  2542 => x"c84a717c",
  2543 => x"48722ab7",
  2544 => x"7098ffc3",
  2545 => x"d04a717c",
  2546 => x"48722ab7",
  2547 => x"7098ffc3",
  2548 => x"d848717c",
  2549 => x"7c7028b7",
  2550 => x"7c7c7cc0",
  2551 => x"7c7c7c7c",
  2552 => x"7c7c7c7c",
  2553 => x"48d0ff7c",
  2554 => x"c478e0c0",
  2555 => x"49dc1e66",
  2556 => x"87d1d8ff",
  2557 => x"8efc86c8",
  2558 => x"4c264d26",
  2559 => x"4f264b26",
  2560 => x"d0e0c21e",
  2561 => x"defe49bf",
  2562 => x"48c087c0",
  2563 => x"00004f26",
  2564 => x"00002814",
  2565 => x"32434956",
  2566 => x"20202030",
  2567 => x"004d4f52",
  2568 => x"00001bb3",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
