
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"f3",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"dc",x"f3",x"c2"),
    18 => (x"48",x"e4",x"e0",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"e4",x"e0",x"c2",x"87"),
    25 => (x"e0",x"e0",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e8",x"c1",x"87",x"f7"),
    29 => (x"e0",x"c2",x"87",x"ca"),
    30 => (x"e0",x"c2",x"4d",x"e4"),
    31 => (x"ad",x"74",x"4c",x"e4"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"d0",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"c3",x"4c",x"87",x"ca"),
    69 => (x"74",x"9c",x"98",x"df"),
    70 => (x"87",x"eb",x"02",x"88"),
    71 => (x"4b",x"26",x"4a",x"26"),
    72 => (x"4f",x"26",x"4c",x"26"),
    73 => (x"81",x"48",x"73",x"1e"),
    74 => (x"c5",x"02",x"a9",x"73"),
    75 => (x"05",x"53",x"12",x"87"),
    76 => (x"4f",x"26",x"87",x"f6"),
    77 => (x"71",x"1e",x"73",x"1e"),
    78 => (x"4b",x"66",x"c8",x"4a"),
    79 => (x"71",x"8b",x"c1",x"49"),
    80 => (x"87",x"cf",x"02",x"99"),
    81 => (x"d4",x"ff",x"48",x"12"),
    82 => (x"49",x"73",x"78",x"08"),
    83 => (x"99",x"71",x"8b",x"c1"),
    84 => (x"26",x"87",x"f1",x"05"),
    85 => (x"0e",x"4f",x"26",x"4b"),
    86 => (x"0e",x"5c",x"5b",x"5e"),
    87 => (x"d4",x"ff",x"4a",x"71"),
    88 => (x"4b",x"66",x"cc",x"4c"),
    89 => (x"71",x"8b",x"c1",x"49"),
    90 => (x"87",x"ce",x"02",x"99"),
    91 => (x"6c",x"7c",x"ff",x"c3"),
    92 => (x"c1",x"49",x"73",x"52"),
    93 => (x"05",x"99",x"71",x"8b"),
    94 => (x"4c",x"26",x"87",x"f2"),
    95 => (x"4f",x"26",x"4b",x"26"),
    96 => (x"ff",x"1e",x"73",x"1e"),
    97 => (x"ff",x"c3",x"4b",x"d4"),
    98 => (x"c3",x"4a",x"6b",x"7b"),
    99 => (x"49",x"6b",x"7b",x"ff"),
   100 => (x"b1",x"72",x"32",x"c8"),
   101 => (x"6b",x"7b",x"ff",x"c3"),
   102 => (x"71",x"31",x"c8",x"4a"),
   103 => (x"7b",x"ff",x"c3",x"b2"),
   104 => (x"32",x"c8",x"49",x"6b"),
   105 => (x"48",x"71",x"b1",x"72"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4d",x"71",x"0e",x"5d"),
   109 => (x"75",x"4c",x"d4",x"ff"),
   110 => (x"98",x"ff",x"c3",x"48"),
   111 => (x"e0",x"c2",x"7c",x"70"),
   112 => (x"c8",x"05",x"bf",x"e4"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"48",x"71",x"29",x"d8"),
   117 => (x"70",x"98",x"ff",x"c3"),
   118 => (x"49",x"66",x"d0",x"7c"),
   119 => (x"48",x"71",x"29",x"d0"),
   120 => (x"70",x"98",x"ff",x"c3"),
   121 => (x"49",x"66",x"d0",x"7c"),
   122 => (x"48",x"71",x"29",x"c8"),
   123 => (x"70",x"98",x"ff",x"c3"),
   124 => (x"48",x"66",x"d0",x"7c"),
   125 => (x"70",x"98",x"ff",x"c3"),
   126 => (x"d0",x"49",x"75",x"7c"),
   127 => (x"c3",x"48",x"71",x"29"),
   128 => (x"7c",x"70",x"98",x"ff"),
   129 => (x"f0",x"c9",x"4b",x"6c"),
   130 => (x"ff",x"c3",x"4a",x"ff"),
   131 => (x"87",x"cf",x"05",x"ab"),
   132 => (x"6c",x"7c",x"71",x"49"),
   133 => (x"02",x"8a",x"c1",x"4b"),
   134 => (x"ab",x"71",x"87",x"c5"),
   135 => (x"73",x"87",x"f2",x"02"),
   136 => (x"26",x"4d",x"26",x"48"),
   137 => (x"26",x"4b",x"26",x"4c"),
   138 => (x"49",x"c0",x"1e",x"4f"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"81",x"c1",x"78",x"ff"),
   141 => (x"a9",x"b7",x"c8",x"c3"),
   142 => (x"26",x"87",x"f1",x"04"),
   143 => (x"5b",x"5e",x"0e",x"4f"),
   144 => (x"c0",x"0e",x"5d",x"5c"),
   145 => (x"f7",x"c1",x"f0",x"ff"),
   146 => (x"c0",x"c0",x"c1",x"4d"),
   147 => (x"4b",x"c0",x"c0",x"c0"),
   148 => (x"c4",x"87",x"d6",x"ff"),
   149 => (x"c0",x"4c",x"df",x"f8"),
   150 => (x"fd",x"49",x"75",x"1e"),
   151 => (x"86",x"c4",x"87",x"ce"),
   152 => (x"c0",x"05",x"a8",x"c1"),
   153 => (x"d4",x"ff",x"87",x"e5"),
   154 => (x"78",x"ff",x"c3",x"48"),
   155 => (x"e1",x"c0",x"1e",x"73"),
   156 => (x"49",x"e9",x"c1",x"f0"),
   157 => (x"c4",x"87",x"f5",x"fc"),
   158 => (x"05",x"98",x"70",x"86"),
   159 => (x"d4",x"ff",x"87",x"ca"),
   160 => (x"78",x"ff",x"c3",x"48"),
   161 => (x"87",x"cb",x"48",x"c1"),
   162 => (x"c1",x"87",x"de",x"fe"),
   163 => (x"c6",x"ff",x"05",x"8c"),
   164 => (x"26",x"48",x"c0",x"87"),
   165 => (x"26",x"4c",x"26",x"4d"),
   166 => (x"0e",x"4f",x"26",x"4b"),
   167 => (x"0e",x"5c",x"5b",x"5e"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"d4",x"ff",x"4c",x"c1"),
   170 => (x"78",x"ff",x"c3",x"48"),
   171 => (x"f7",x"49",x"e0",x"cb"),
   172 => (x"4b",x"d3",x"87",x"f5"),
   173 => (x"49",x"74",x"1e",x"c0"),
   174 => (x"c4",x"87",x"f1",x"fb"),
   175 => (x"05",x"98",x"70",x"86"),
   176 => (x"d4",x"ff",x"87",x"ca"),
   177 => (x"78",x"ff",x"c3",x"48"),
   178 => (x"87",x"cb",x"48",x"c1"),
   179 => (x"c1",x"87",x"da",x"fd"),
   180 => (x"df",x"ff",x"05",x"8b"),
   181 => (x"26",x"48",x"c0",x"87"),
   182 => (x"26",x"4b",x"26",x"4c"),
   183 => (x"00",x"00",x"00",x"4f"),
   184 => (x"00",x"44",x"4d",x"43"),
   185 => (x"5c",x"5b",x"5e",x"0e"),
   186 => (x"ff",x"c3",x"0e",x"5d"),
   187 => (x"4b",x"d4",x"ff",x"4d"),
   188 => (x"c6",x"87",x"f6",x"fc"),
   189 => (x"e1",x"c0",x"1e",x"ea"),
   190 => (x"49",x"c8",x"c1",x"f0"),
   191 => (x"c4",x"87",x"ed",x"fa"),
   192 => (x"02",x"a8",x"c1",x"86"),
   193 => (x"d2",x"fe",x"87",x"c8"),
   194 => (x"c1",x"48",x"c0",x"87"),
   195 => (x"ef",x"f9",x"87",x"e8"),
   196 => (x"cf",x"49",x"70",x"87"),
   197 => (x"c6",x"99",x"ff",x"ff"),
   198 => (x"c8",x"02",x"a9",x"ea"),
   199 => (x"87",x"fb",x"fd",x"87"),
   200 => (x"d1",x"c1",x"48",x"c0"),
   201 => (x"c0",x"7b",x"75",x"87"),
   202 => (x"d0",x"fc",x"4c",x"f1"),
   203 => (x"02",x"98",x"70",x"87"),
   204 => (x"c0",x"87",x"ec",x"c0"),
   205 => (x"f0",x"ff",x"c0",x"1e"),
   206 => (x"f9",x"49",x"fa",x"c1"),
   207 => (x"86",x"c4",x"87",x"ee"),
   208 => (x"da",x"05",x"98",x"70"),
   209 => (x"6b",x"7b",x"75",x"87"),
   210 => (x"75",x"7b",x"75",x"49"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"99",x"c0",x"c1",x"7b"),
   213 => (x"c1",x"87",x"c4",x"02"),
   214 => (x"c0",x"87",x"db",x"48"),
   215 => (x"c2",x"87",x"d7",x"48"),
   216 => (x"87",x"ca",x"05",x"ac"),
   217 => (x"f4",x"49",x"c0",x"ce"),
   218 => (x"48",x"c0",x"87",x"fd"),
   219 => (x"8c",x"c1",x"87",x"c8"),
   220 => (x"87",x"f6",x"fe",x"05"),
   221 => (x"4d",x"26",x"48",x"c0"),
   222 => (x"4b",x"26",x"4c",x"26"),
   223 => (x"00",x"00",x"4f",x"26"),
   224 => (x"43",x"48",x"44",x"53"),
   225 => (x"69",x"61",x"66",x"20"),
   226 => (x"00",x"0a",x"21",x"6c"),
   227 => (x"5c",x"5b",x"5e",x"0e"),
   228 => (x"d0",x"ff",x"0e",x"5d"),
   229 => (x"d0",x"e5",x"c0",x"4d"),
   230 => (x"c2",x"4c",x"c0",x"c1"),
   231 => (x"c1",x"48",x"e4",x"e0"),
   232 => (x"49",x"d8",x"d0",x"78"),
   233 => (x"c7",x"87",x"c0",x"f4"),
   234 => (x"f9",x"7d",x"c2",x"4b"),
   235 => (x"7d",x"c3",x"87",x"fb"),
   236 => (x"49",x"74",x"1e",x"c0"),
   237 => (x"c4",x"87",x"f5",x"f7"),
   238 => (x"05",x"a8",x"c1",x"86"),
   239 => (x"c2",x"4b",x"87",x"c1"),
   240 => (x"87",x"cb",x"05",x"ab"),
   241 => (x"f3",x"49",x"d0",x"d0"),
   242 => (x"48",x"c0",x"87",x"dd"),
   243 => (x"c1",x"87",x"f6",x"c0"),
   244 => (x"d4",x"ff",x"05",x"8b"),
   245 => (x"87",x"cc",x"fc",x"87"),
   246 => (x"58",x"e8",x"e0",x"c2"),
   247 => (x"cd",x"05",x"98",x"70"),
   248 => (x"c0",x"1e",x"c1",x"87"),
   249 => (x"d0",x"c1",x"f0",x"ff"),
   250 => (x"87",x"c0",x"f7",x"49"),
   251 => (x"d4",x"ff",x"86",x"c4"),
   252 => (x"78",x"ff",x"c3",x"48"),
   253 => (x"c2",x"87",x"cc",x"c5"),
   254 => (x"c2",x"58",x"ec",x"e0"),
   255 => (x"48",x"d4",x"ff",x"7d"),
   256 => (x"c1",x"78",x"ff",x"c3"),
   257 => (x"26",x"4d",x"26",x"48"),
   258 => (x"26",x"4b",x"26",x"4c"),
   259 => (x"00",x"00",x"00",x"4f"),
   260 => (x"52",x"52",x"45",x"49"),
   261 => (x"00",x"00",x"00",x"00"),
   262 => (x"00",x"49",x"50",x"53"),
   263 => (x"5c",x"5b",x"5e",x"0e"),
   264 => (x"4d",x"71",x"0e",x"5d"),
   265 => (x"ff",x"4c",x"ff",x"c3"),
   266 => (x"7b",x"74",x"4b",x"d4"),
   267 => (x"c4",x"48",x"d0",x"ff"),
   268 => (x"7b",x"74",x"78",x"c3"),
   269 => (x"ff",x"c0",x"1e",x"75"),
   270 => (x"49",x"d8",x"c1",x"f0"),
   271 => (x"c4",x"87",x"ed",x"f5"),
   272 => (x"02",x"98",x"70",x"86"),
   273 => (x"c8",x"d2",x"87",x"cb"),
   274 => (x"87",x"db",x"f1",x"49"),
   275 => (x"ee",x"c0",x"48",x"c1"),
   276 => (x"c3",x"7b",x"74",x"87"),
   277 => (x"c0",x"c8",x"7b",x"fe"),
   278 => (x"49",x"66",x"d4",x"1e"),
   279 => (x"c4",x"87",x"d5",x"f3"),
   280 => (x"74",x"7b",x"74",x"86"),
   281 => (x"d8",x"7b",x"74",x"7b"),
   282 => (x"74",x"4a",x"e0",x"da"),
   283 => (x"c5",x"05",x"6b",x"7b"),
   284 => (x"05",x"8a",x"c1",x"87"),
   285 => (x"7b",x"74",x"87",x"f5"),
   286 => (x"c2",x"48",x"d0",x"ff"),
   287 => (x"26",x"48",x"c0",x"78"),
   288 => (x"26",x"4c",x"26",x"4d"),
   289 => (x"00",x"4f",x"26",x"4b"),
   290 => (x"74",x"69",x"72",x"57"),
   291 => (x"61",x"66",x"20",x"65"),
   292 => (x"64",x"65",x"6c",x"69"),
   293 => (x"5e",x"0e",x"00",x"0a"),
   294 => (x"0e",x"5d",x"5c",x"5b"),
   295 => (x"4b",x"71",x"86",x"fc"),
   296 => (x"c0",x"4c",x"d4",x"ff"),
   297 => (x"cd",x"ee",x"c5",x"7e"),
   298 => (x"ff",x"c3",x"4a",x"df"),
   299 => (x"c3",x"48",x"6c",x"7c"),
   300 => (x"c0",x"05",x"a8",x"fe"),
   301 => (x"4d",x"74",x"87",x"f8"),
   302 => (x"cc",x"02",x"9b",x"73"),
   303 => (x"1e",x"66",x"d4",x"87"),
   304 => (x"d2",x"f2",x"49",x"73"),
   305 => (x"d4",x"86",x"c4",x"87"),
   306 => (x"48",x"d0",x"ff",x"87"),
   307 => (x"d4",x"78",x"d1",x"c4"),
   308 => (x"ff",x"c3",x"4a",x"66"),
   309 => (x"05",x"8a",x"c1",x"7d"),
   310 => (x"a6",x"d8",x"87",x"f8"),
   311 => (x"7c",x"ff",x"c3",x"5a"),
   312 => (x"05",x"9b",x"73",x"7c"),
   313 => (x"d0",x"ff",x"87",x"c5"),
   314 => (x"c1",x"78",x"d0",x"48"),
   315 => (x"8a",x"c1",x"7e",x"4a"),
   316 => (x"87",x"f6",x"fe",x"05"),
   317 => (x"8e",x"fc",x"48",x"6e"),
   318 => (x"4c",x"26",x"4d",x"26"),
   319 => (x"4f",x"26",x"4b",x"26"),
   320 => (x"71",x"1e",x"73",x"1e"),
   321 => (x"ff",x"4b",x"c0",x"4a"),
   322 => (x"ff",x"c3",x"48",x"d4"),
   323 => (x"48",x"d0",x"ff",x"78"),
   324 => (x"ff",x"78",x"c3",x"c4"),
   325 => (x"ff",x"c3",x"48",x"d4"),
   326 => (x"c0",x"1e",x"72",x"78"),
   327 => (x"d1",x"c1",x"f0",x"ff"),
   328 => (x"87",x"c8",x"f2",x"49"),
   329 => (x"98",x"70",x"86",x"c4"),
   330 => (x"c8",x"87",x"d2",x"05"),
   331 => (x"66",x"cc",x"1e",x"c0"),
   332 => (x"87",x"e2",x"fd",x"49"),
   333 => (x"4b",x"70",x"86",x"c4"),
   334 => (x"c2",x"48",x"d0",x"ff"),
   335 => (x"26",x"48",x"73",x"78"),
   336 => (x"0e",x"4f",x"26",x"4b"),
   337 => (x"5d",x"5c",x"5b",x"5e"),
   338 => (x"c0",x"1e",x"c0",x"0e"),
   339 => (x"c9",x"c1",x"f0",x"ff"),
   340 => (x"87",x"d8",x"f1",x"49"),
   341 => (x"e0",x"c2",x"1e",x"d2"),
   342 => (x"f9",x"fc",x"49",x"ec"),
   343 => (x"c0",x"86",x"c8",x"87"),
   344 => (x"d2",x"84",x"c1",x"4c"),
   345 => (x"f8",x"04",x"ac",x"b7"),
   346 => (x"ec",x"e0",x"c2",x"87"),
   347 => (x"c3",x"49",x"bf",x"97"),
   348 => (x"c0",x"c1",x"99",x"c0"),
   349 => (x"e7",x"c0",x"05",x"a9"),
   350 => (x"f3",x"e0",x"c2",x"87"),
   351 => (x"d0",x"49",x"bf",x"97"),
   352 => (x"f4",x"e0",x"c2",x"31"),
   353 => (x"c8",x"4a",x"bf",x"97"),
   354 => (x"c2",x"b1",x"72",x"32"),
   355 => (x"bf",x"97",x"f5",x"e0"),
   356 => (x"4c",x"71",x"b1",x"4a"),
   357 => (x"ff",x"ff",x"ff",x"cf"),
   358 => (x"ca",x"84",x"c1",x"9c"),
   359 => (x"87",x"e7",x"c1",x"34"),
   360 => (x"97",x"f5",x"e0",x"c2"),
   361 => (x"31",x"c1",x"49",x"bf"),
   362 => (x"e0",x"c2",x"99",x"c6"),
   363 => (x"4a",x"bf",x"97",x"f6"),
   364 => (x"72",x"2a",x"b7",x"c7"),
   365 => (x"f1",x"e0",x"c2",x"b1"),
   366 => (x"4d",x"4a",x"bf",x"97"),
   367 => (x"e0",x"c2",x"9d",x"cf"),
   368 => (x"4a",x"bf",x"97",x"f2"),
   369 => (x"32",x"ca",x"9a",x"c3"),
   370 => (x"97",x"f3",x"e0",x"c2"),
   371 => (x"33",x"c2",x"4b",x"bf"),
   372 => (x"e0",x"c2",x"b2",x"73"),
   373 => (x"4b",x"bf",x"97",x"f4"),
   374 => (x"c6",x"9b",x"c0",x"c3"),
   375 => (x"b2",x"73",x"2b",x"b7"),
   376 => (x"48",x"c1",x"81",x"c2"),
   377 => (x"49",x"70",x"30",x"71"),
   378 => (x"30",x"75",x"48",x"c1"),
   379 => (x"4c",x"72",x"4d",x"70"),
   380 => (x"94",x"71",x"84",x"c1"),
   381 => (x"ad",x"b7",x"c0",x"c8"),
   382 => (x"c1",x"87",x"cc",x"06"),
   383 => (x"c8",x"2d",x"b7",x"34"),
   384 => (x"01",x"ad",x"b7",x"c0"),
   385 => (x"74",x"87",x"f4",x"ff"),
   386 => (x"26",x"4d",x"26",x"48"),
   387 => (x"26",x"4b",x"26",x"4c"),
   388 => (x"5b",x"5e",x"0e",x"4f"),
   389 => (x"f8",x"0e",x"5d",x"5c"),
   390 => (x"d4",x"e9",x"c2",x"86"),
   391 => (x"c2",x"78",x"c0",x"48"),
   392 => (x"c0",x"1e",x"cc",x"e1"),
   393 => (x"87",x"d8",x"fb",x"49"),
   394 => (x"98",x"70",x"86",x"c4"),
   395 => (x"c0",x"87",x"c5",x"05"),
   396 => (x"87",x"c0",x"c9",x"48"),
   397 => (x"7e",x"c1",x"4d",x"c0"),
   398 => (x"bf",x"dc",x"f7",x"c0"),
   399 => (x"c2",x"e2",x"c2",x"49"),
   400 => (x"4b",x"c8",x"71",x"4a"),
   401 => (x"70",x"87",x"df",x"ea"),
   402 => (x"87",x"c2",x"05",x"98"),
   403 => (x"f7",x"c0",x"7e",x"c0"),
   404 => (x"c2",x"49",x"bf",x"d8"),
   405 => (x"71",x"4a",x"de",x"e2"),
   406 => (x"c9",x"ea",x"4b",x"c8"),
   407 => (x"05",x"98",x"70",x"87"),
   408 => (x"7e",x"c0",x"87",x"c2"),
   409 => (x"fd",x"c0",x"02",x"6e"),
   410 => (x"d2",x"e8",x"c2",x"87"),
   411 => (x"e9",x"c2",x"4d",x"bf"),
   412 => (x"7e",x"bf",x"9f",x"ca"),
   413 => (x"ea",x"d6",x"c5",x"48"),
   414 => (x"87",x"c7",x"05",x"a8"),
   415 => (x"bf",x"d2",x"e8",x"c2"),
   416 => (x"6e",x"87",x"ce",x"4d"),
   417 => (x"d5",x"e9",x"ca",x"48"),
   418 => (x"87",x"c5",x"02",x"a8"),
   419 => (x"e3",x"c7",x"48",x"c0"),
   420 => (x"cc",x"e1",x"c2",x"87"),
   421 => (x"f9",x"49",x"75",x"1e"),
   422 => (x"86",x"c4",x"87",x"e6"),
   423 => (x"c5",x"05",x"98",x"70"),
   424 => (x"c7",x"48",x"c0",x"87"),
   425 => (x"f7",x"c0",x"87",x"ce"),
   426 => (x"c2",x"49",x"bf",x"d8"),
   427 => (x"71",x"4a",x"de",x"e2"),
   428 => (x"f1",x"e8",x"4b",x"c8"),
   429 => (x"05",x"98",x"70",x"87"),
   430 => (x"e9",x"c2",x"87",x"c8"),
   431 => (x"78",x"c1",x"48",x"d4"),
   432 => (x"f7",x"c0",x"87",x"da"),
   433 => (x"c2",x"49",x"bf",x"dc"),
   434 => (x"71",x"4a",x"c2",x"e2"),
   435 => (x"d5",x"e8",x"4b",x"c8"),
   436 => (x"02",x"98",x"70",x"87"),
   437 => (x"c0",x"87",x"c5",x"c0"),
   438 => (x"87",x"d8",x"c6",x"48"),
   439 => (x"97",x"ca",x"e9",x"c2"),
   440 => (x"d5",x"c1",x"49",x"bf"),
   441 => (x"cd",x"c0",x"05",x"a9"),
   442 => (x"cb",x"e9",x"c2",x"87"),
   443 => (x"c2",x"49",x"bf",x"97"),
   444 => (x"c0",x"02",x"a9",x"ea"),
   445 => (x"48",x"c0",x"87",x"c5"),
   446 => (x"c2",x"87",x"f9",x"c5"),
   447 => (x"bf",x"97",x"cc",x"e1"),
   448 => (x"e9",x"c3",x"48",x"7e"),
   449 => (x"ce",x"c0",x"02",x"a8"),
   450 => (x"c3",x"48",x"6e",x"87"),
   451 => (x"c0",x"02",x"a8",x"eb"),
   452 => (x"48",x"c0",x"87",x"c5"),
   453 => (x"c2",x"87",x"dd",x"c5"),
   454 => (x"bf",x"97",x"d7",x"e1"),
   455 => (x"c0",x"05",x"99",x"49"),
   456 => (x"e1",x"c2",x"87",x"cc"),
   457 => (x"49",x"bf",x"97",x"d8"),
   458 => (x"c0",x"02",x"a9",x"c2"),
   459 => (x"48",x"c0",x"87",x"c5"),
   460 => (x"c2",x"87",x"c1",x"c5"),
   461 => (x"bf",x"97",x"d9",x"e1"),
   462 => (x"d0",x"e9",x"c2",x"48"),
   463 => (x"48",x"4c",x"70",x"58"),
   464 => (x"e9",x"c2",x"88",x"c1"),
   465 => (x"e1",x"c2",x"58",x"d4"),
   466 => (x"49",x"bf",x"97",x"da"),
   467 => (x"e1",x"c2",x"81",x"75"),
   468 => (x"4a",x"bf",x"97",x"db"),
   469 => (x"a1",x"72",x"32",x"c8"),
   470 => (x"e4",x"ed",x"c2",x"7e"),
   471 => (x"c2",x"78",x"6e",x"48"),
   472 => (x"bf",x"97",x"dc",x"e1"),
   473 => (x"58",x"a6",x"c8",x"48"),
   474 => (x"bf",x"d4",x"e9",x"c2"),
   475 => (x"87",x"cf",x"c2",x"02"),
   476 => (x"bf",x"d8",x"f7",x"c0"),
   477 => (x"de",x"e2",x"c2",x"49"),
   478 => (x"4b",x"c8",x"71",x"4a"),
   479 => (x"70",x"87",x"e7",x"e5"),
   480 => (x"c5",x"c0",x"02",x"98"),
   481 => (x"c3",x"48",x"c0",x"87"),
   482 => (x"e9",x"c2",x"87",x"ea"),
   483 => (x"c2",x"4c",x"bf",x"cc"),
   484 => (x"c2",x"5c",x"f8",x"ed"),
   485 => (x"bf",x"97",x"f1",x"e1"),
   486 => (x"c2",x"31",x"c8",x"49"),
   487 => (x"bf",x"97",x"f0",x"e1"),
   488 => (x"c2",x"49",x"a1",x"4a"),
   489 => (x"bf",x"97",x"f2",x"e1"),
   490 => (x"72",x"32",x"d0",x"4a"),
   491 => (x"e1",x"c2",x"49",x"a1"),
   492 => (x"4a",x"bf",x"97",x"f3"),
   493 => (x"a1",x"72",x"32",x"d8"),
   494 => (x"91",x"66",x"c4",x"49"),
   495 => (x"bf",x"e4",x"ed",x"c2"),
   496 => (x"ec",x"ed",x"c2",x"81"),
   497 => (x"f9",x"e1",x"c2",x"59"),
   498 => (x"c8",x"4a",x"bf",x"97"),
   499 => (x"f8",x"e1",x"c2",x"32"),
   500 => (x"a2",x"4b",x"bf",x"97"),
   501 => (x"fa",x"e1",x"c2",x"4a"),
   502 => (x"d0",x"4b",x"bf",x"97"),
   503 => (x"4a",x"a2",x"73",x"33"),
   504 => (x"97",x"fb",x"e1",x"c2"),
   505 => (x"9b",x"cf",x"4b",x"bf"),
   506 => (x"a2",x"73",x"33",x"d8"),
   507 => (x"f0",x"ed",x"c2",x"4a"),
   508 => (x"74",x"8a",x"c2",x"5a"),
   509 => (x"f0",x"ed",x"c2",x"92"),
   510 => (x"78",x"a1",x"72",x"48"),
   511 => (x"c2",x"87",x"c1",x"c1"),
   512 => (x"bf",x"97",x"de",x"e1"),
   513 => (x"c2",x"31",x"c8",x"49"),
   514 => (x"bf",x"97",x"dd",x"e1"),
   515 => (x"c5",x"49",x"a1",x"4a"),
   516 => (x"81",x"ff",x"c7",x"31"),
   517 => (x"ed",x"c2",x"29",x"c9"),
   518 => (x"e1",x"c2",x"59",x"f8"),
   519 => (x"4a",x"bf",x"97",x"e3"),
   520 => (x"e1",x"c2",x"32",x"c8"),
   521 => (x"4b",x"bf",x"97",x"e2"),
   522 => (x"66",x"c4",x"4a",x"a2"),
   523 => (x"c2",x"82",x"6e",x"92"),
   524 => (x"c2",x"5a",x"f4",x"ed"),
   525 => (x"c0",x"48",x"ec",x"ed"),
   526 => (x"e8",x"ed",x"c2",x"78"),
   527 => (x"78",x"a1",x"72",x"48"),
   528 => (x"48",x"f8",x"ed",x"c2"),
   529 => (x"bf",x"ec",x"ed",x"c2"),
   530 => (x"fc",x"ed",x"c2",x"78"),
   531 => (x"f0",x"ed",x"c2",x"48"),
   532 => (x"e9",x"c2",x"78",x"bf"),
   533 => (x"c0",x"02",x"bf",x"d4"),
   534 => (x"48",x"74",x"87",x"c9"),
   535 => (x"7e",x"70",x"30",x"c4"),
   536 => (x"c2",x"87",x"c9",x"c0"),
   537 => (x"48",x"bf",x"f4",x"ed"),
   538 => (x"7e",x"70",x"30",x"c4"),
   539 => (x"48",x"d8",x"e9",x"c2"),
   540 => (x"48",x"c1",x"78",x"6e"),
   541 => (x"4d",x"26",x"8e",x"f8"),
   542 => (x"4b",x"26",x"4c",x"26"),
   543 => (x"5e",x"0e",x"4f",x"26"),
   544 => (x"0e",x"5d",x"5c",x"5b"),
   545 => (x"e9",x"c2",x"4a",x"71"),
   546 => (x"cb",x"02",x"bf",x"d4"),
   547 => (x"c7",x"4b",x"72",x"87"),
   548 => (x"c1",x"4d",x"72",x"2b"),
   549 => (x"87",x"c9",x"9d",x"ff"),
   550 => (x"2b",x"c8",x"4b",x"72"),
   551 => (x"ff",x"c3",x"4d",x"72"),
   552 => (x"e4",x"ed",x"c2",x"9d"),
   553 => (x"f7",x"c0",x"83",x"bf"),
   554 => (x"02",x"ab",x"bf",x"d4"),
   555 => (x"f7",x"c0",x"87",x"d9"),
   556 => (x"e1",x"c2",x"5b",x"d8"),
   557 => (x"49",x"73",x"1e",x"cc"),
   558 => (x"c4",x"87",x"c5",x"f1"),
   559 => (x"05",x"98",x"70",x"86"),
   560 => (x"48",x"c0",x"87",x"c5"),
   561 => (x"c2",x"87",x"e6",x"c0"),
   562 => (x"02",x"bf",x"d4",x"e9"),
   563 => (x"49",x"75",x"87",x"d2"),
   564 => (x"e1",x"c2",x"91",x"c4"),
   565 => (x"4c",x"69",x"81",x"cc"),
   566 => (x"ff",x"ff",x"ff",x"cf"),
   567 => (x"87",x"cb",x"9c",x"ff"),
   568 => (x"91",x"c2",x"49",x"75"),
   569 => (x"81",x"cc",x"e1",x"c2"),
   570 => (x"74",x"4c",x"69",x"9f"),
   571 => (x"26",x"4d",x"26",x"48"),
   572 => (x"26",x"4b",x"26",x"4c"),
   573 => (x"5b",x"5e",x"0e",x"4f"),
   574 => (x"f4",x"0e",x"5d",x"5c"),
   575 => (x"59",x"a6",x"cc",x"86"),
   576 => (x"c5",x"05",x"66",x"c8"),
   577 => (x"c3",x"48",x"c0",x"87"),
   578 => (x"66",x"c8",x"87",x"c8"),
   579 => (x"70",x"80",x"c8",x"48"),
   580 => (x"78",x"c0",x"48",x"7e"),
   581 => (x"c7",x"02",x"66",x"dc"),
   582 => (x"97",x"66",x"dc",x"87"),
   583 => (x"87",x"c5",x"05",x"bf"),
   584 => (x"ed",x"c2",x"48",x"c0"),
   585 => (x"c1",x"1e",x"c0",x"87"),
   586 => (x"ee",x"ca",x"49",x"49"),
   587 => (x"70",x"86",x"c4",x"87"),
   588 => (x"c0",x"02",x"9c",x"4c"),
   589 => (x"e9",x"c2",x"87",x"fc"),
   590 => (x"66",x"dc",x"4a",x"dc"),
   591 => (x"ca",x"de",x"ff",x"49"),
   592 => (x"02",x"98",x"70",x"87"),
   593 => (x"74",x"87",x"eb",x"c0"),
   594 => (x"49",x"66",x"dc",x"4a"),
   595 => (x"de",x"ff",x"4b",x"cb"),
   596 => (x"98",x"70",x"87",x"ee"),
   597 => (x"c0",x"87",x"db",x"02"),
   598 => (x"02",x"9c",x"74",x"1e"),
   599 => (x"4d",x"c0",x"87",x"c4"),
   600 => (x"4d",x"c1",x"87",x"c2"),
   601 => (x"f2",x"c9",x"49",x"75"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"ff",x"05",x"9c",x"4c"),
   604 => (x"9c",x"74",x"87",x"c4"),
   605 => (x"87",x"d8",x"c1",x"02"),
   606 => (x"6e",x"49",x"a4",x"dc"),
   607 => (x"da",x"78",x"69",x"48"),
   608 => (x"66",x"c8",x"49",x"a4"),
   609 => (x"c8",x"80",x"c4",x"48"),
   610 => (x"69",x"9f",x"58",x"a6"),
   611 => (x"08",x"66",x"c4",x"48"),
   612 => (x"d4",x"e9",x"c2",x"78"),
   613 => (x"87",x"d2",x"02",x"bf"),
   614 => (x"9f",x"49",x"a4",x"d4"),
   615 => (x"ff",x"c0",x"49",x"69"),
   616 => (x"48",x"71",x"99",x"ff"),
   617 => (x"7e",x"70",x"30",x"d0"),
   618 => (x"7e",x"c0",x"87",x"c2"),
   619 => (x"c4",x"48",x"49",x"6e"),
   620 => (x"c4",x"80",x"bf",x"66"),
   621 => (x"c8",x"78",x"08",x"66"),
   622 => (x"78",x"c0",x"48",x"66"),
   623 => (x"cc",x"49",x"66",x"c8"),
   624 => (x"bf",x"66",x"c4",x"81"),
   625 => (x"49",x"66",x"c8",x"79"),
   626 => (x"79",x"c0",x"81",x"d0"),
   627 => (x"87",x"c2",x"48",x"c1"),
   628 => (x"8e",x"f4",x"48",x"c0"),
   629 => (x"4c",x"26",x"4d",x"26"),
   630 => (x"4f",x"26",x"4b",x"26"),
   631 => (x"5c",x"5b",x"5e",x"0e"),
   632 => (x"4c",x"71",x"0e",x"5d"),
   633 => (x"74",x"4d",x"66",x"d0"),
   634 => (x"c6",x"c1",x"02",x"9c"),
   635 => (x"49",x"a4",x"c8",x"87"),
   636 => (x"fe",x"c0",x"02",x"69"),
   637 => (x"6c",x"4a",x"75",x"87"),
   638 => (x"4d",x"a1",x"72",x"49"),
   639 => (x"d0",x"e9",x"c2",x"b9"),
   640 => (x"ba",x"ff",x"4a",x"bf"),
   641 => (x"99",x"71",x"99",x"72"),
   642 => (x"87",x"e5",x"c0",x"02"),
   643 => (x"6b",x"4b",x"a4",x"c4"),
   644 => (x"87",x"ea",x"f9",x"49"),
   645 => (x"e9",x"c2",x"7b",x"70"),
   646 => (x"6c",x"49",x"bf",x"cc"),
   647 => (x"75",x"7c",x"71",x"81"),
   648 => (x"e9",x"c2",x"b9",x"4a"),
   649 => (x"ff",x"4a",x"bf",x"d0"),
   650 => (x"71",x"99",x"72",x"ba"),
   651 => (x"db",x"ff",x"05",x"99"),
   652 => (x"26",x"7c",x"75",x"87"),
   653 => (x"26",x"4c",x"26",x"4d"),
   654 => (x"1e",x"4f",x"26",x"4b"),
   655 => (x"4b",x"71",x"1e",x"73"),
   656 => (x"87",x"c7",x"02",x"9b"),
   657 => (x"69",x"49",x"a3",x"c8"),
   658 => (x"c0",x"87",x"c5",x"05"),
   659 => (x"87",x"f6",x"c0",x"48"),
   660 => (x"bf",x"e8",x"ed",x"c2"),
   661 => (x"4a",x"a3",x"c4",x"49"),
   662 => (x"8a",x"c2",x"4a",x"6a"),
   663 => (x"bf",x"cc",x"e9",x"c2"),
   664 => (x"49",x"a1",x"72",x"92"),
   665 => (x"bf",x"d0",x"e9",x"c2"),
   666 => (x"72",x"9a",x"6b",x"4a"),
   667 => (x"f7",x"c0",x"49",x"a1"),
   668 => (x"66",x"c8",x"59",x"d8"),
   669 => (x"c7",x"ea",x"71",x"1e"),
   670 => (x"70",x"86",x"c4",x"87"),
   671 => (x"87",x"c4",x"05",x"98"),
   672 => (x"87",x"c2",x"48",x"c0"),
   673 => (x"4b",x"26",x"48",x"c1"),
   674 => (x"73",x"1e",x"4f",x"26"),
   675 => (x"9b",x"4b",x"71",x"1e"),
   676 => (x"c8",x"87",x"c7",x"02"),
   677 => (x"05",x"69",x"49",x"a3"),
   678 => (x"48",x"c0",x"87",x"c5"),
   679 => (x"c2",x"87",x"f6",x"c0"),
   680 => (x"49",x"bf",x"e8",x"ed"),
   681 => (x"6a",x"4a",x"a3",x"c4"),
   682 => (x"c2",x"8a",x"c2",x"4a"),
   683 => (x"92",x"bf",x"cc",x"e9"),
   684 => (x"c2",x"49",x"a1",x"72"),
   685 => (x"4a",x"bf",x"d0",x"e9"),
   686 => (x"a1",x"72",x"9a",x"6b"),
   687 => (x"d8",x"f7",x"c0",x"49"),
   688 => (x"1e",x"66",x"c8",x"59"),
   689 => (x"87",x"d4",x"e5",x"71"),
   690 => (x"98",x"70",x"86",x"c4"),
   691 => (x"c0",x"87",x"c4",x"05"),
   692 => (x"c1",x"87",x"c2",x"48"),
   693 => (x"26",x"4b",x"26",x"48"),
   694 => (x"5b",x"5e",x"0e",x"4f"),
   695 => (x"fc",x"0e",x"5d",x"5c"),
   696 => (x"d4",x"4b",x"71",x"86"),
   697 => (x"9b",x"73",x"4d",x"66"),
   698 => (x"87",x"cc",x"c1",x"02"),
   699 => (x"69",x"49",x"a3",x"c8"),
   700 => (x"87",x"c4",x"c1",x"02"),
   701 => (x"c2",x"4c",x"a3",x"d0"),
   702 => (x"49",x"bf",x"d0",x"e9"),
   703 => (x"4a",x"6c",x"b9",x"ff"),
   704 => (x"66",x"d4",x"7e",x"99"),
   705 => (x"87",x"cd",x"06",x"a9"),
   706 => (x"cc",x"7c",x"7b",x"c0"),
   707 => (x"a3",x"c4",x"4a",x"a3"),
   708 => (x"ca",x"79",x"6a",x"49"),
   709 => (x"f8",x"49",x"72",x"87"),
   710 => (x"66",x"d4",x"99",x"c0"),
   711 => (x"75",x"8d",x"71",x"4d"),
   712 => (x"71",x"29",x"c9",x"49"),
   713 => (x"fa",x"49",x"73",x"1e"),
   714 => (x"e1",x"c2",x"87",x"f2"),
   715 => (x"49",x"73",x"1e",x"cc"),
   716 => (x"c8",x"87",x"c8",x"fc"),
   717 => (x"7c",x"66",x"d4",x"86"),
   718 => (x"4d",x"26",x"8e",x"fc"),
   719 => (x"4b",x"26",x"4c",x"26"),
   720 => (x"73",x"1e",x"4f",x"26"),
   721 => (x"9b",x"4b",x"71",x"1e"),
   722 => (x"87",x"e4",x"c0",x"02"),
   723 => (x"5b",x"fc",x"ed",x"c2"),
   724 => (x"8a",x"c2",x"4a",x"73"),
   725 => (x"bf",x"cc",x"e9",x"c2"),
   726 => (x"ed",x"c2",x"92",x"49"),
   727 => (x"72",x"48",x"bf",x"e8"),
   728 => (x"c0",x"ee",x"c2",x"80"),
   729 => (x"c4",x"48",x"71",x"58"),
   730 => (x"dc",x"e9",x"c2",x"30"),
   731 => (x"87",x"ed",x"c0",x"58"),
   732 => (x"48",x"f8",x"ed",x"c2"),
   733 => (x"bf",x"ec",x"ed",x"c2"),
   734 => (x"fc",x"ed",x"c2",x"78"),
   735 => (x"f0",x"ed",x"c2",x"48"),
   736 => (x"e9",x"c2",x"78",x"bf"),
   737 => (x"c9",x"02",x"bf",x"d4"),
   738 => (x"cc",x"e9",x"c2",x"87"),
   739 => (x"31",x"c4",x"49",x"bf"),
   740 => (x"ed",x"c2",x"87",x"c7"),
   741 => (x"c4",x"49",x"bf",x"f4"),
   742 => (x"dc",x"e9",x"c2",x"31"),
   743 => (x"26",x"4b",x"26",x"59"),
   744 => (x"5b",x"5e",x"0e",x"4f"),
   745 => (x"4a",x"71",x"0e",x"5c"),
   746 => (x"9a",x"72",x"4b",x"c0"),
   747 => (x"87",x"e0",x"c0",x"02"),
   748 => (x"9f",x"49",x"a2",x"da"),
   749 => (x"e9",x"c2",x"4b",x"69"),
   750 => (x"cf",x"02",x"bf",x"d4"),
   751 => (x"49",x"a2",x"d4",x"87"),
   752 => (x"4c",x"49",x"69",x"9f"),
   753 => (x"9c",x"ff",x"ff",x"c0"),
   754 => (x"87",x"c2",x"34",x"d0"),
   755 => (x"b3",x"74",x"4c",x"c0"),
   756 => (x"ed",x"fd",x"49",x"73"),
   757 => (x"26",x"4c",x"26",x"87"),
   758 => (x"0e",x"4f",x"26",x"4b"),
   759 => (x"5d",x"5c",x"5b",x"5e"),
   760 => (x"c8",x"86",x"f0",x"0e"),
   761 => (x"ff",x"cf",x"59",x"a6"),
   762 => (x"4c",x"f8",x"ff",x"ff"),
   763 => (x"66",x"c4",x"7e",x"c0"),
   764 => (x"c2",x"87",x"d8",x"02"),
   765 => (x"c0",x"48",x"c8",x"e1"),
   766 => (x"c0",x"e1",x"c2",x"78"),
   767 => (x"fc",x"ed",x"c2",x"48"),
   768 => (x"e1",x"c2",x"78",x"bf"),
   769 => (x"ed",x"c2",x"48",x"c4"),
   770 => (x"c2",x"78",x"bf",x"f8"),
   771 => (x"c0",x"48",x"e9",x"e9"),
   772 => (x"d8",x"e9",x"c2",x"50"),
   773 => (x"e1",x"c2",x"49",x"bf"),
   774 => (x"71",x"4a",x"bf",x"c8"),
   775 => (x"cb",x"c4",x"03",x"aa"),
   776 => (x"cf",x"49",x"72",x"87"),
   777 => (x"e9",x"c0",x"05",x"99"),
   778 => (x"d4",x"f7",x"c0",x"87"),
   779 => (x"c0",x"e1",x"c2",x"48"),
   780 => (x"e1",x"c2",x"78",x"bf"),
   781 => (x"e1",x"c2",x"1e",x"cc"),
   782 => (x"c2",x"49",x"bf",x"c0"),
   783 => (x"c1",x"48",x"c0",x"e1"),
   784 => (x"e2",x"71",x"78",x"a1"),
   785 => (x"86",x"c4",x"87",x"fa"),
   786 => (x"48",x"d0",x"f7",x"c0"),
   787 => (x"78",x"cc",x"e1",x"c2"),
   788 => (x"f7",x"c0",x"87",x"cc"),
   789 => (x"c0",x"48",x"bf",x"d0"),
   790 => (x"f7",x"c0",x"80",x"e0"),
   791 => (x"e1",x"c2",x"58",x"d4"),
   792 => (x"c1",x"48",x"bf",x"c8"),
   793 => (x"cc",x"e1",x"c2",x"80"),
   794 => (x"0d",x"d0",x"27",x"58"),
   795 => (x"97",x"bf",x"00",x"00"),
   796 => (x"02",x"9d",x"4d",x"bf"),
   797 => (x"c3",x"87",x"e5",x"c2"),
   798 => (x"c2",x"02",x"ad",x"e5"),
   799 => (x"f7",x"c0",x"87",x"de"),
   800 => (x"cb",x"4b",x"bf",x"d0"),
   801 => (x"4c",x"11",x"49",x"a3"),
   802 => (x"c1",x"05",x"ac",x"cf"),
   803 => (x"49",x"75",x"87",x"d2"),
   804 => (x"89",x"c1",x"99",x"df"),
   805 => (x"e9",x"c2",x"91",x"cd"),
   806 => (x"a3",x"c1",x"81",x"dc"),
   807 => (x"c3",x"51",x"12",x"4a"),
   808 => (x"51",x"12",x"4a",x"a3"),
   809 => (x"12",x"4a",x"a3",x"c5"),
   810 => (x"4a",x"a3",x"c7",x"51"),
   811 => (x"a3",x"c9",x"51",x"12"),
   812 => (x"ce",x"51",x"12",x"4a"),
   813 => (x"51",x"12",x"4a",x"a3"),
   814 => (x"12",x"4a",x"a3",x"d0"),
   815 => (x"4a",x"a3",x"d2",x"51"),
   816 => (x"a3",x"d4",x"51",x"12"),
   817 => (x"d6",x"51",x"12",x"4a"),
   818 => (x"51",x"12",x"4a",x"a3"),
   819 => (x"12",x"4a",x"a3",x"d8"),
   820 => (x"4a",x"a3",x"dc",x"51"),
   821 => (x"a3",x"de",x"51",x"12"),
   822 => (x"c1",x"51",x"12",x"4a"),
   823 => (x"87",x"fc",x"c0",x"7e"),
   824 => (x"99",x"c8",x"49",x"74"),
   825 => (x"87",x"ed",x"c0",x"05"),
   826 => (x"99",x"d0",x"49",x"74"),
   827 => (x"c0",x"87",x"d3",x"05"),
   828 => (x"c0",x"02",x"66",x"e0"),
   829 => (x"49",x"73",x"87",x"cc"),
   830 => (x"0f",x"66",x"e0",x"c0"),
   831 => (x"c0",x"02",x"98",x"70"),
   832 => (x"05",x"6e",x"87",x"d3"),
   833 => (x"c2",x"87",x"c6",x"c0"),
   834 => (x"c0",x"48",x"dc",x"e9"),
   835 => (x"d0",x"f7",x"c0",x"50"),
   836 => (x"eb",x"c2",x"48",x"bf"),
   837 => (x"e9",x"e9",x"c2",x"87"),
   838 => (x"7e",x"50",x"c0",x"48"),
   839 => (x"bf",x"d8",x"e9",x"c2"),
   840 => (x"c8",x"e1",x"c2",x"49"),
   841 => (x"aa",x"71",x"4a",x"bf"),
   842 => (x"87",x"f5",x"fb",x"04"),
   843 => (x"ff",x"ff",x"ff",x"cf"),
   844 => (x"ed",x"c2",x"4c",x"f8"),
   845 => (x"c0",x"05",x"bf",x"fc"),
   846 => (x"e9",x"c2",x"87",x"c8"),
   847 => (x"c1",x"02",x"bf",x"d4"),
   848 => (x"e1",x"c2",x"87",x"fc"),
   849 => (x"ec",x"49",x"bf",x"c4"),
   850 => (x"e1",x"c2",x"87",x"f4"),
   851 => (x"a6",x"c4",x"58",x"c8"),
   852 => (x"c4",x"e1",x"c2",x"48"),
   853 => (x"e9",x"c2",x"78",x"bf"),
   854 => (x"c0",x"02",x"bf",x"d4"),
   855 => (x"66",x"c4",x"87",x"db"),
   856 => (x"74",x"99",x"74",x"49"),
   857 => (x"c8",x"c0",x"02",x"a9"),
   858 => (x"48",x"a6",x"c8",x"87"),
   859 => (x"e7",x"c0",x"78",x"c0"),
   860 => (x"48",x"a6",x"c8",x"87"),
   861 => (x"df",x"c0",x"78",x"c1"),
   862 => (x"49",x"66",x"c4",x"87"),
   863 => (x"99",x"f8",x"ff",x"cf"),
   864 => (x"c8",x"c0",x"02",x"a9"),
   865 => (x"48",x"a6",x"cc",x"87"),
   866 => (x"c5",x"c0",x"78",x"c0"),
   867 => (x"48",x"a6",x"cc",x"87"),
   868 => (x"a6",x"c8",x"78",x"c1"),
   869 => (x"78",x"66",x"cc",x"48"),
   870 => (x"c0",x"05",x"66",x"c8"),
   871 => (x"66",x"c4",x"87",x"e0"),
   872 => (x"c2",x"89",x"c2",x"49"),
   873 => (x"4a",x"bf",x"cc",x"e9"),
   874 => (x"e8",x"ed",x"c2",x"91"),
   875 => (x"e1",x"c2",x"4a",x"bf"),
   876 => (x"a1",x"72",x"48",x"c0"),
   877 => (x"c8",x"e1",x"c2",x"78"),
   878 => (x"f9",x"78",x"c0",x"48"),
   879 => (x"48",x"c0",x"87",x"d3"),
   880 => (x"ff",x"ff",x"ff",x"cf"),
   881 => (x"8e",x"f0",x"4c",x"f8"),
   882 => (x"4c",x"26",x"4d",x"26"),
   883 => (x"4f",x"26",x"4b",x"26"),
   884 => (x"00",x"00",x"00",x"00"),
   885 => (x"ff",x"ff",x"ff",x"ff"),
   886 => (x"00",x"00",x"0d",x"e0"),
   887 => (x"00",x"00",x"0d",x"ec"),
   888 => (x"33",x"54",x"41",x"46"),
   889 => (x"20",x"20",x"20",x"32"),
   890 => (x"00",x"00",x"00",x"00"),
   891 => (x"31",x"54",x"41",x"46"),
   892 => (x"20",x"20",x"20",x"36"),
   893 => (x"d4",x"ff",x"1e",x"00"),
   894 => (x"78",x"ff",x"c3",x"48"),
   895 => (x"4f",x"26",x"48",x"68"),
   896 => (x"48",x"d4",x"ff",x"1e"),
   897 => (x"ff",x"78",x"ff",x"c3"),
   898 => (x"e1",x"c0",x"48",x"d0"),
   899 => (x"48",x"d4",x"ff",x"78"),
   900 => (x"4f",x"26",x"78",x"d4"),
   901 => (x"48",x"d0",x"ff",x"1e"),
   902 => (x"26",x"78",x"e0",x"c0"),
   903 => (x"d4",x"ff",x"1e",x"4f"),
   904 => (x"99",x"49",x"70",x"87"),
   905 => (x"c0",x"87",x"c6",x"02"),
   906 => (x"f1",x"05",x"a9",x"fb"),
   907 => (x"26",x"48",x"71",x"87"),
   908 => (x"5b",x"5e",x"0e",x"4f"),
   909 => (x"4b",x"71",x"0e",x"5c"),
   910 => (x"f8",x"fe",x"4c",x"c0"),
   911 => (x"99",x"49",x"70",x"87"),
   912 => (x"87",x"f9",x"c0",x"02"),
   913 => (x"02",x"a9",x"ec",x"c0"),
   914 => (x"c0",x"87",x"f2",x"c0"),
   915 => (x"c0",x"02",x"a9",x"fb"),
   916 => (x"66",x"cc",x"87",x"eb"),
   917 => (x"c7",x"03",x"ac",x"b7"),
   918 => (x"02",x"66",x"d0",x"87"),
   919 => (x"53",x"71",x"87",x"c2"),
   920 => (x"c2",x"02",x"99",x"71"),
   921 => (x"fe",x"84",x"c1",x"87"),
   922 => (x"49",x"70",x"87",x"cb"),
   923 => (x"87",x"cd",x"02",x"99"),
   924 => (x"02",x"a9",x"ec",x"c0"),
   925 => (x"fb",x"c0",x"87",x"c7"),
   926 => (x"d5",x"ff",x"05",x"a9"),
   927 => (x"02",x"66",x"d0",x"87"),
   928 => (x"97",x"c0",x"87",x"c3"),
   929 => (x"a9",x"ec",x"c0",x"7b"),
   930 => (x"74",x"87",x"c4",x"05"),
   931 => (x"74",x"87",x"c5",x"4a"),
   932 => (x"8a",x"0a",x"c0",x"4a"),
   933 => (x"4c",x"26",x"48",x"72"),
   934 => (x"4f",x"26",x"4b",x"26"),
   935 => (x"87",x"d5",x"fd",x"1e"),
   936 => (x"c0",x"4a",x"49",x"70"),
   937 => (x"c9",x"04",x"aa",x"f0"),
   938 => (x"aa",x"f9",x"c0",x"87"),
   939 => (x"c0",x"87",x"c3",x"01"),
   940 => (x"c1",x"c1",x"8a",x"f0"),
   941 => (x"87",x"c9",x"04",x"aa"),
   942 => (x"01",x"aa",x"da",x"c1"),
   943 => (x"f7",x"c0",x"87",x"c3"),
   944 => (x"26",x"48",x"72",x"8a"),
   945 => (x"5b",x"5e",x"0e",x"4f"),
   946 => (x"f8",x"0e",x"5d",x"5c"),
   947 => (x"c0",x"4c",x"71",x"86"),
   948 => (x"87",x"ec",x"fc",x"7e"),
   949 => (x"fd",x"c0",x"4b",x"c0"),
   950 => (x"49",x"bf",x"97",x"e4"),
   951 => (x"cf",x"04",x"a9",x"c0"),
   952 => (x"87",x"f9",x"fc",x"87"),
   953 => (x"fd",x"c0",x"83",x"c1"),
   954 => (x"49",x"bf",x"97",x"e4"),
   955 => (x"87",x"f1",x"06",x"ab"),
   956 => (x"97",x"e4",x"fd",x"c0"),
   957 => (x"87",x"cf",x"02",x"bf"),
   958 => (x"70",x"87",x"fa",x"fb"),
   959 => (x"c6",x"02",x"99",x"49"),
   960 => (x"a9",x"ec",x"c0",x"87"),
   961 => (x"c0",x"87",x"f1",x"05"),
   962 => (x"87",x"e9",x"fb",x"4b"),
   963 => (x"e4",x"fb",x"4d",x"70"),
   964 => (x"58",x"a6",x"c8",x"87"),
   965 => (x"70",x"87",x"de",x"fb"),
   966 => (x"c8",x"83",x"c1",x"4a"),
   967 => (x"69",x"97",x"49",x"a4"),
   968 => (x"da",x"05",x"ad",x"49"),
   969 => (x"49",x"a4",x"c9",x"87"),
   970 => (x"c4",x"49",x"69",x"97"),
   971 => (x"ce",x"05",x"a9",x"66"),
   972 => (x"49",x"a4",x"ca",x"87"),
   973 => (x"aa",x"49",x"69",x"97"),
   974 => (x"c1",x"87",x"c4",x"05"),
   975 => (x"c0",x"87",x"d0",x"7e"),
   976 => (x"c6",x"02",x"ad",x"ec"),
   977 => (x"ad",x"fb",x"c0",x"87"),
   978 => (x"c0",x"87",x"c4",x"05"),
   979 => (x"6e",x"7e",x"c1",x"4b"),
   980 => (x"87",x"f5",x"fe",x"02"),
   981 => (x"73",x"87",x"fd",x"fa"),
   982 => (x"26",x"8e",x"f8",x"48"),
   983 => (x"26",x"4c",x"26",x"4d"),
   984 => (x"00",x"4f",x"26",x"4b"),
   985 => (x"1e",x"73",x"1e",x"00"),
   986 => (x"c8",x"4b",x"d4",x"ff"),
   987 => (x"d0",x"ff",x"4a",x"66"),
   988 => (x"78",x"c5",x"c8",x"48"),
   989 => (x"c1",x"48",x"d4",x"ff"),
   990 => (x"7b",x"11",x"78",x"d4"),
   991 => (x"f9",x"05",x"8a",x"c1"),
   992 => (x"48",x"d0",x"ff",x"87"),
   993 => (x"4b",x"26",x"78",x"c4"),
   994 => (x"5e",x"0e",x"4f",x"26"),
   995 => (x"0e",x"5d",x"5c",x"5b"),
   996 => (x"7e",x"71",x"86",x"f8"),
   997 => (x"ee",x"c2",x"1e",x"6e"),
   998 => (x"d8",x"e5",x"49",x"cc"),
   999 => (x"70",x"86",x"c4",x"87"),
  1000 => (x"e4",x"c4",x"02",x"98"),
  1001 => (x"ec",x"ec",x"c1",x"87"),
  1002 => (x"49",x"6e",x"4c",x"bf"),
  1003 => (x"c8",x"87",x"d6",x"fc"),
  1004 => (x"98",x"70",x"58",x"a6"),
  1005 => (x"c4",x"87",x"c5",x"05"),
  1006 => (x"78",x"c1",x"48",x"a6"),
  1007 => (x"c5",x"48",x"d0",x"ff"),
  1008 => (x"48",x"d4",x"ff",x"78"),
  1009 => (x"c4",x"78",x"d5",x"c1"),
  1010 => (x"89",x"c1",x"49",x"66"),
  1011 => (x"ec",x"c1",x"31",x"c6"),
  1012 => (x"4a",x"bf",x"97",x"e4"),
  1013 => (x"ff",x"b0",x"71",x"48"),
  1014 => (x"ff",x"78",x"08",x"d4"),
  1015 => (x"78",x"c4",x"48",x"d0"),
  1016 => (x"97",x"c8",x"ee",x"c2"),
  1017 => (x"99",x"d0",x"49",x"bf"),
  1018 => (x"c5",x"87",x"dd",x"02"),
  1019 => (x"48",x"d4",x"ff",x"78"),
  1020 => (x"c0",x"78",x"d6",x"c1"),
  1021 => (x"48",x"d4",x"ff",x"4a"),
  1022 => (x"c1",x"78",x"ff",x"c3"),
  1023 => (x"aa",x"e0",x"c0",x"82"),
  1024 => (x"ff",x"87",x"f2",x"04"),
  1025 => (x"78",x"c4",x"48",x"d0"),
  1026 => (x"c3",x"48",x"d4",x"ff"),
  1027 => (x"d0",x"ff",x"78",x"ff"),
  1028 => (x"ff",x"78",x"c5",x"48"),
  1029 => (x"d3",x"c1",x"48",x"d4"),
  1030 => (x"ff",x"78",x"c1",x"78"),
  1031 => (x"78",x"c4",x"48",x"d0"),
  1032 => (x"06",x"ac",x"b7",x"c0"),
  1033 => (x"c2",x"87",x"cb",x"c2"),
  1034 => (x"4b",x"bf",x"d4",x"ee"),
  1035 => (x"73",x"7e",x"74",x"8c"),
  1036 => (x"dd",x"c1",x"02",x"9b"),
  1037 => (x"4d",x"c0",x"c8",x"87"),
  1038 => (x"ab",x"b7",x"c0",x"8b"),
  1039 => (x"c8",x"87",x"c6",x"03"),
  1040 => (x"c0",x"4d",x"a3",x"c0"),
  1041 => (x"c8",x"ee",x"c2",x"4b"),
  1042 => (x"d0",x"49",x"bf",x"97"),
  1043 => (x"87",x"cf",x"02",x"99"),
  1044 => (x"ee",x"c2",x"1e",x"c0"),
  1045 => (x"e2",x"e7",x"49",x"cc"),
  1046 => (x"70",x"86",x"c4",x"87"),
  1047 => (x"c2",x"87",x"d8",x"4c"),
  1048 => (x"c2",x"1e",x"cc",x"e1"),
  1049 => (x"e7",x"49",x"cc",x"ee"),
  1050 => (x"4c",x"70",x"87",x"d1"),
  1051 => (x"e1",x"c2",x"1e",x"75"),
  1052 => (x"f0",x"fb",x"49",x"cc"),
  1053 => (x"74",x"86",x"c8",x"87"),
  1054 => (x"87",x"c5",x"05",x"9c"),
  1055 => (x"ca",x"c1",x"48",x"c0"),
  1056 => (x"c2",x"1e",x"c1",x"87"),
  1057 => (x"e5",x"49",x"cc",x"ee"),
  1058 => (x"86",x"c4",x"87",x"d2"),
  1059 => (x"fe",x"05",x"9b",x"73"),
  1060 => (x"4c",x"6e",x"87",x"e3"),
  1061 => (x"06",x"ac",x"b7",x"c0"),
  1062 => (x"ee",x"c2",x"87",x"d1"),
  1063 => (x"78",x"c0",x"48",x"cc"),
  1064 => (x"78",x"c0",x"80",x"d0"),
  1065 => (x"ee",x"c2",x"80",x"f4"),
  1066 => (x"c0",x"78",x"bf",x"d8"),
  1067 => (x"fd",x"01",x"ac",x"b7"),
  1068 => (x"d0",x"ff",x"87",x"f5"),
  1069 => (x"ff",x"78",x"c5",x"48"),
  1070 => (x"d3",x"c1",x"48",x"d4"),
  1071 => (x"ff",x"78",x"c0",x"78"),
  1072 => (x"78",x"c4",x"48",x"d0"),
  1073 => (x"c2",x"c0",x"48",x"c1"),
  1074 => (x"f8",x"48",x"c0",x"87"),
  1075 => (x"26",x"4d",x"26",x"8e"),
  1076 => (x"26",x"4b",x"26",x"4c"),
  1077 => (x"5b",x"5e",x"0e",x"4f"),
  1078 => (x"fc",x"0e",x"5d",x"5c"),
  1079 => (x"c0",x"4d",x"71",x"86"),
  1080 => (x"04",x"ad",x"4c",x"4b"),
  1081 => (x"c0",x"87",x"e8",x"c0"),
  1082 => (x"74",x"1e",x"c5",x"fb"),
  1083 => (x"87",x"c4",x"02",x"9c"),
  1084 => (x"87",x"c2",x"4a",x"c0"),
  1085 => (x"49",x"72",x"4a",x"c1"),
  1086 => (x"c4",x"87",x"e0",x"eb"),
  1087 => (x"c1",x"7e",x"70",x"86"),
  1088 => (x"c2",x"05",x"6e",x"83"),
  1089 => (x"c1",x"4b",x"75",x"87"),
  1090 => (x"06",x"ab",x"75",x"84"),
  1091 => (x"6e",x"87",x"d8",x"ff"),
  1092 => (x"26",x"8e",x"fc",x"48"),
  1093 => (x"26",x"4c",x"26",x"4d"),
  1094 => (x"0e",x"4f",x"26",x"4b"),
  1095 => (x"0e",x"5c",x"5b",x"5e"),
  1096 => (x"66",x"cc",x"4b",x"71"),
  1097 => (x"4c",x"87",x"d8",x"02"),
  1098 => (x"02",x"8c",x"f0",x"c0"),
  1099 => (x"4a",x"74",x"87",x"d8"),
  1100 => (x"d1",x"02",x"8a",x"c1"),
  1101 => (x"cd",x"02",x"8a",x"87"),
  1102 => (x"c9",x"02",x"8a",x"87"),
  1103 => (x"73",x"87",x"d9",x"87"),
  1104 => (x"87",x"c6",x"f9",x"49"),
  1105 => (x"1e",x"74",x"87",x"d2"),
  1106 => (x"d8",x"c1",x"49",x"c0"),
  1107 => (x"1e",x"74",x"87",x"ee"),
  1108 => (x"d8",x"c1",x"49",x"73"),
  1109 => (x"86",x"c8",x"87",x"e6"),
  1110 => (x"4b",x"26",x"4c",x"26"),
  1111 => (x"5e",x"0e",x"4f",x"26"),
  1112 => (x"0e",x"5d",x"5c",x"5b"),
  1113 => (x"4c",x"71",x"86",x"fc"),
  1114 => (x"c2",x"91",x"de",x"49"),
  1115 => (x"71",x"4d",x"f8",x"ee"),
  1116 => (x"02",x"6d",x"97",x"85"),
  1117 => (x"c2",x"87",x"dc",x"c1"),
  1118 => (x"49",x"bf",x"e8",x"ee"),
  1119 => (x"fd",x"71",x"81",x"74"),
  1120 => (x"7e",x"70",x"87",x"d3"),
  1121 => (x"c0",x"02",x"98",x"48"),
  1122 => (x"ee",x"c2",x"87",x"f2"),
  1123 => (x"4a",x"70",x"4b",x"ec"),
  1124 => (x"fe",x"fe",x"49",x"cb"),
  1125 => (x"4b",x"74",x"87",x"ce"),
  1126 => (x"ec",x"c1",x"93",x"cc"),
  1127 => (x"83",x"c4",x"83",x"f0"),
  1128 => (x"7b",x"e0",x"c7",x"c1"),
  1129 => (x"c3",x"c1",x"49",x"74"),
  1130 => (x"7b",x"75",x"87",x"de"),
  1131 => (x"97",x"e8",x"ec",x"c1"),
  1132 => (x"c2",x"1e",x"49",x"bf"),
  1133 => (x"fd",x"49",x"ec",x"ee"),
  1134 => (x"86",x"c4",x"87",x"e1"),
  1135 => (x"c3",x"c1",x"49",x"74"),
  1136 => (x"49",x"c0",x"87",x"c6"),
  1137 => (x"87",x"e1",x"c4",x"c1"),
  1138 => (x"48",x"c4",x"ee",x"c2"),
  1139 => (x"c0",x"49",x"50",x"c0"),
  1140 => (x"fc",x"87",x"cc",x"e2"),
  1141 => (x"26",x"4d",x"26",x"8e"),
  1142 => (x"26",x"4b",x"26",x"4c"),
  1143 => (x"00",x"00",x"00",x"4f"),
  1144 => (x"64",x"61",x"6f",x"4c"),
  1145 => (x"2e",x"67",x"6e",x"69"),
  1146 => (x"1e",x"00",x"2e",x"2e"),
  1147 => (x"4b",x"71",x"1e",x"73"),
  1148 => (x"e8",x"ee",x"c2",x"49"),
  1149 => (x"fb",x"71",x"81",x"bf"),
  1150 => (x"4a",x"70",x"87",x"db"),
  1151 => (x"87",x"c4",x"02",x"9a"),
  1152 => (x"87",x"dd",x"e6",x"49"),
  1153 => (x"48",x"e8",x"ee",x"c2"),
  1154 => (x"49",x"73",x"78",x"c0"),
  1155 => (x"26",x"87",x"fa",x"c1"),
  1156 => (x"1e",x"4f",x"26",x"4b"),
  1157 => (x"4b",x"71",x"1e",x"73"),
  1158 => (x"02",x"4a",x"a3",x"c4"),
  1159 => (x"c1",x"87",x"d0",x"c1"),
  1160 => (x"87",x"dc",x"02",x"8a"),
  1161 => (x"f2",x"c0",x"02",x"8a"),
  1162 => (x"c1",x"05",x"8a",x"87"),
  1163 => (x"ee",x"c2",x"87",x"d3"),
  1164 => (x"c1",x"02",x"bf",x"e8"),
  1165 => (x"c1",x"48",x"87",x"cb"),
  1166 => (x"ec",x"ee",x"c2",x"88"),
  1167 => (x"87",x"c1",x"c1",x"58"),
  1168 => (x"bf",x"e8",x"ee",x"c2"),
  1169 => (x"c2",x"89",x"c6",x"49"),
  1170 => (x"c0",x"59",x"ec",x"ee"),
  1171 => (x"c0",x"03",x"a9",x"b7"),
  1172 => (x"ee",x"c2",x"87",x"ef"),
  1173 => (x"78",x"c0",x"48",x"e8"),
  1174 => (x"c2",x"87",x"e6",x"c0"),
  1175 => (x"02",x"bf",x"e4",x"ee"),
  1176 => (x"ee",x"c2",x"87",x"df"),
  1177 => (x"c1",x"48",x"bf",x"e8"),
  1178 => (x"ec",x"ee",x"c2",x"80"),
  1179 => (x"c2",x"87",x"d2",x"58"),
  1180 => (x"02",x"bf",x"e4",x"ee"),
  1181 => (x"ee",x"c2",x"87",x"cb"),
  1182 => (x"c6",x"48",x"bf",x"e8"),
  1183 => (x"ec",x"ee",x"c2",x"80"),
  1184 => (x"c4",x"49",x"73",x"58"),
  1185 => (x"26",x"4b",x"26",x"87"),
  1186 => (x"5b",x"5e",x"0e",x"4f"),
  1187 => (x"f0",x"0e",x"5d",x"5c"),
  1188 => (x"59",x"a6",x"d0",x"86"),
  1189 => (x"4d",x"cc",x"e1",x"c2"),
  1190 => (x"ee",x"c2",x"4c",x"c0"),
  1191 => (x"78",x"c1",x"48",x"e4"),
  1192 => (x"c0",x"48",x"a6",x"c4"),
  1193 => (x"c2",x"7e",x"75",x"78"),
  1194 => (x"48",x"bf",x"e8",x"ee"),
  1195 => (x"c0",x"06",x"a8",x"c0"),
  1196 => (x"7e",x"75",x"87",x"fa"),
  1197 => (x"48",x"cc",x"e1",x"c2"),
  1198 => (x"ef",x"c0",x"02",x"98"),
  1199 => (x"c5",x"fb",x"c0",x"87"),
  1200 => (x"02",x"66",x"c8",x"1e"),
  1201 => (x"4d",x"c0",x"87",x"c4"),
  1202 => (x"4d",x"c1",x"87",x"c2"),
  1203 => (x"ca",x"e4",x"49",x"75"),
  1204 => (x"70",x"86",x"c4",x"87"),
  1205 => (x"c4",x"84",x"c1",x"7e"),
  1206 => (x"80",x"c1",x"48",x"66"),
  1207 => (x"c2",x"58",x"a6",x"c8"),
  1208 => (x"ac",x"bf",x"e8",x"ee"),
  1209 => (x"6e",x"87",x"c5",x"03"),
  1210 => (x"87",x"d1",x"ff",x"05"),
  1211 => (x"4c",x"c0",x"4d",x"6e"),
  1212 => (x"c3",x"02",x"9d",x"75"),
  1213 => (x"fb",x"c0",x"87",x"e0"),
  1214 => (x"66",x"c8",x"1e",x"c5"),
  1215 => (x"cc",x"87",x"c7",x"02"),
  1216 => (x"78",x"c0",x"48",x"a6"),
  1217 => (x"a6",x"cc",x"87",x"c5"),
  1218 => (x"cc",x"78",x"c1",x"48"),
  1219 => (x"ca",x"e3",x"49",x"66"),
  1220 => (x"70",x"86",x"c4",x"87"),
  1221 => (x"02",x"98",x"48",x"7e"),
  1222 => (x"49",x"87",x"e8",x"c2"),
  1223 => (x"69",x"97",x"81",x"cb"),
  1224 => (x"02",x"99",x"d0",x"49"),
  1225 => (x"c1",x"87",x"d6",x"c1"),
  1226 => (x"74",x"4a",x"eb",x"c7"),
  1227 => (x"c1",x"91",x"cc",x"49"),
  1228 => (x"72",x"81",x"f0",x"ec"),
  1229 => (x"c3",x"81",x"c8",x"79"),
  1230 => (x"49",x"74",x"51",x"ff"),
  1231 => (x"ee",x"c2",x"91",x"de"),
  1232 => (x"85",x"71",x"4d",x"f8"),
  1233 => (x"7d",x"97",x"c1",x"c2"),
  1234 => (x"c0",x"49",x"a5",x"c1"),
  1235 => (x"e9",x"c2",x"51",x"e0"),
  1236 => (x"02",x"bf",x"97",x"dc"),
  1237 => (x"84",x"c1",x"87",x"d2"),
  1238 => (x"c2",x"4b",x"a5",x"c2"),
  1239 => (x"db",x"4a",x"dc",x"e9"),
  1240 => (x"ff",x"f6",x"fe",x"49"),
  1241 => (x"87",x"db",x"c1",x"87"),
  1242 => (x"c0",x"49",x"a5",x"cd"),
  1243 => (x"c2",x"84",x"c1",x"51"),
  1244 => (x"4a",x"6e",x"4b",x"a5"),
  1245 => (x"f6",x"fe",x"49",x"cb"),
  1246 => (x"c6",x"c1",x"87",x"ea"),
  1247 => (x"de",x"c5",x"c1",x"87"),
  1248 => (x"cc",x"49",x"74",x"4a"),
  1249 => (x"f0",x"ec",x"c1",x"91"),
  1250 => (x"c2",x"79",x"72",x"81"),
  1251 => (x"bf",x"97",x"dc",x"e9"),
  1252 => (x"74",x"87",x"d8",x"02"),
  1253 => (x"c1",x"91",x"de",x"49"),
  1254 => (x"f8",x"ee",x"c2",x"84"),
  1255 => (x"c2",x"83",x"71",x"4b"),
  1256 => (x"dd",x"4a",x"dc",x"e9"),
  1257 => (x"fb",x"f5",x"fe",x"49"),
  1258 => (x"74",x"87",x"d8",x"87"),
  1259 => (x"c2",x"93",x"de",x"4b"),
  1260 => (x"cb",x"83",x"f8",x"ee"),
  1261 => (x"51",x"c0",x"49",x"a3"),
  1262 => (x"6e",x"73",x"84",x"c1"),
  1263 => (x"fe",x"49",x"cb",x"4a"),
  1264 => (x"c4",x"87",x"e1",x"f5"),
  1265 => (x"80",x"c1",x"48",x"66"),
  1266 => (x"c7",x"58",x"a6",x"c8"),
  1267 => (x"c5",x"c0",x"03",x"ac"),
  1268 => (x"fc",x"05",x"6e",x"87"),
  1269 => (x"ac",x"c7",x"87",x"e0"),
  1270 => (x"87",x"e6",x"c0",x"03"),
  1271 => (x"48",x"e4",x"ee",x"c2"),
  1272 => (x"c5",x"c1",x"78",x"c0"),
  1273 => (x"49",x"74",x"4a",x"de"),
  1274 => (x"ec",x"c1",x"91",x"cc"),
  1275 => (x"79",x"72",x"81",x"f0"),
  1276 => (x"91",x"de",x"49",x"74"),
  1277 => (x"81",x"f8",x"ee",x"c2"),
  1278 => (x"84",x"c1",x"51",x"c0"),
  1279 => (x"ff",x"04",x"ac",x"c7"),
  1280 => (x"ee",x"c1",x"87",x"da"),
  1281 => (x"50",x"c0",x"48",x"cc"),
  1282 => (x"d1",x"c1",x"80",x"f7"),
  1283 => (x"d0",x"c1",x"40",x"f9"),
  1284 => (x"80",x"c8",x"78",x"ec"),
  1285 => (x"78",x"d3",x"c8",x"c1"),
  1286 => (x"c0",x"49",x"66",x"cc"),
  1287 => (x"f0",x"87",x"e9",x"f9"),
  1288 => (x"26",x"4d",x"26",x"8e"),
  1289 => (x"26",x"4b",x"26",x"4c"),
  1290 => (x"00",x"00",x"00",x"4f"),
  1291 => (x"61",x"42",x"20",x"80"),
  1292 => (x"1e",x"00",x"6b",x"63"),
  1293 => (x"4b",x"71",x"1e",x"73"),
  1294 => (x"c1",x"91",x"cc",x"49"),
  1295 => (x"c8",x"81",x"f0",x"ec"),
  1296 => (x"ec",x"c1",x"4a",x"a1"),
  1297 => (x"50",x"12",x"48",x"e4"),
  1298 => (x"c0",x"4a",x"a1",x"c9"),
  1299 => (x"12",x"48",x"e4",x"fd"),
  1300 => (x"c1",x"81",x"ca",x"50"),
  1301 => (x"11",x"48",x"e8",x"ec"),
  1302 => (x"e8",x"ec",x"c1",x"50"),
  1303 => (x"1e",x"49",x"bf",x"97"),
  1304 => (x"f6",x"f2",x"49",x"c0"),
  1305 => (x"f8",x"49",x"73",x"87"),
  1306 => (x"8e",x"fc",x"87",x"df"),
  1307 => (x"4f",x"26",x"4b",x"26"),
  1308 => (x"c0",x"49",x"c0",x"1e"),
  1309 => (x"26",x"87",x"f2",x"f9"),
  1310 => (x"4a",x"71",x"1e",x"4f"),
  1311 => (x"c1",x"91",x"cc",x"49"),
  1312 => (x"c8",x"81",x"f0",x"ec"),
  1313 => (x"c4",x"ee",x"c2",x"81"),
  1314 => (x"c0",x"50",x"11",x"48"),
  1315 => (x"fe",x"49",x"a2",x"f0"),
  1316 => (x"c0",x"87",x"f9",x"ef"),
  1317 => (x"87",x"c7",x"d7",x"49"),
  1318 => (x"ff",x"1e",x"4f",x"26"),
  1319 => (x"ff",x"c3",x"4a",x"d4"),
  1320 => (x"48",x"d0",x"ff",x"7a"),
  1321 => (x"de",x"78",x"e1",x"c0"),
  1322 => (x"48",x"7a",x"71",x"7a"),
  1323 => (x"70",x"28",x"b7",x"c8"),
  1324 => (x"d0",x"48",x"71",x"7a"),
  1325 => (x"7a",x"70",x"28",x"b7"),
  1326 => (x"b7",x"d8",x"48",x"71"),
  1327 => (x"ff",x"7a",x"70",x"28"),
  1328 => (x"e0",x"c0",x"48",x"d0"),
  1329 => (x"0e",x"4f",x"26",x"78"),
  1330 => (x"5d",x"5c",x"5b",x"5e"),
  1331 => (x"71",x"86",x"f4",x"0e"),
  1332 => (x"91",x"cc",x"49",x"4d"),
  1333 => (x"81",x"f0",x"ec",x"c1"),
  1334 => (x"ca",x"4a",x"a1",x"c8"),
  1335 => (x"a6",x"c4",x"7e",x"a1"),
  1336 => (x"c0",x"ee",x"c2",x"48"),
  1337 => (x"97",x"6e",x"78",x"bf"),
  1338 => (x"66",x"c4",x"4b",x"bf"),
  1339 => (x"12",x"2c",x"73",x"4c"),
  1340 => (x"58",x"a6",x"cc",x"48"),
  1341 => (x"84",x"c1",x"9c",x"70"),
  1342 => (x"69",x"97",x"81",x"c9"),
  1343 => (x"04",x"ac",x"b7",x"49"),
  1344 => (x"4c",x"c0",x"87",x"c2"),
  1345 => (x"4a",x"bf",x"97",x"6e"),
  1346 => (x"72",x"49",x"66",x"c8"),
  1347 => (x"c4",x"b9",x"ff",x"31"),
  1348 => (x"48",x"74",x"99",x"66"),
  1349 => (x"4a",x"70",x"30",x"72"),
  1350 => (x"c4",x"ee",x"c2",x"b1"),
  1351 => (x"f9",x"fd",x"71",x"59"),
  1352 => (x"c2",x"1e",x"c7",x"87"),
  1353 => (x"1e",x"bf",x"e0",x"ee"),
  1354 => (x"1e",x"f0",x"ec",x"c1"),
  1355 => (x"97",x"c4",x"ee",x"c2"),
  1356 => (x"f4",x"c1",x"49",x"bf"),
  1357 => (x"c0",x"49",x"75",x"87"),
  1358 => (x"e8",x"87",x"cd",x"f5"),
  1359 => (x"26",x"4d",x"26",x"8e"),
  1360 => (x"26",x"4b",x"26",x"4c"),
  1361 => (x"1e",x"73",x"1e",x"4f"),
  1362 => (x"fd",x"49",x"4b",x"71"),
  1363 => (x"49",x"73",x"87",x"f9"),
  1364 => (x"26",x"87",x"f4",x"fd"),
  1365 => (x"1e",x"4f",x"26",x"4b"),
  1366 => (x"4b",x"71",x"1e",x"73"),
  1367 => (x"02",x"4a",x"a3",x"c2"),
  1368 => (x"8a",x"c1",x"87",x"d6"),
  1369 => (x"87",x"e2",x"c0",x"05"),
  1370 => (x"bf",x"e0",x"ee",x"c2"),
  1371 => (x"48",x"87",x"db",x"02"),
  1372 => (x"ee",x"c2",x"88",x"c1"),
  1373 => (x"87",x"d2",x"58",x"e4"),
  1374 => (x"bf",x"e4",x"ee",x"c2"),
  1375 => (x"c2",x"87",x"cb",x"02"),
  1376 => (x"48",x"bf",x"e0",x"ee"),
  1377 => (x"ee",x"c2",x"80",x"c1"),
  1378 => (x"1e",x"c7",x"58",x"e4"),
  1379 => (x"bf",x"e0",x"ee",x"c2"),
  1380 => (x"f0",x"ec",x"c1",x"1e"),
  1381 => (x"c4",x"ee",x"c2",x"1e"),
  1382 => (x"cc",x"49",x"bf",x"97"),
  1383 => (x"c0",x"49",x"73",x"87"),
  1384 => (x"f4",x"87",x"e5",x"f3"),
  1385 => (x"26",x"4b",x"26",x"8e"),
  1386 => (x"5b",x"5e",x"0e",x"4f"),
  1387 => (x"ff",x"0e",x"5d",x"5c"),
  1388 => (x"e4",x"c0",x"86",x"cc"),
  1389 => (x"a6",x"cc",x"59",x"a6"),
  1390 => (x"c4",x"78",x"c0",x"48"),
  1391 => (x"c4",x"78",x"c0",x"80"),
  1392 => (x"66",x"c8",x"c1",x"80"),
  1393 => (x"c1",x"80",x"c4",x"78"),
  1394 => (x"c1",x"80",x"c4",x"78"),
  1395 => (x"e4",x"ee",x"c2",x"78"),
  1396 => (x"e0",x"78",x"c1",x"48"),
  1397 => (x"c4",x"e1",x"87",x"ea"),
  1398 => (x"87",x"d9",x"e0",x"87"),
  1399 => (x"fb",x"c0",x"4c",x"70"),
  1400 => (x"f3",x"c1",x"02",x"ac"),
  1401 => (x"66",x"e0",x"c0",x"87"),
  1402 => (x"87",x"e8",x"c1",x"05"),
  1403 => (x"4a",x"66",x"c4",x"c1"),
  1404 => (x"7e",x"6a",x"82",x"c4"),
  1405 => (x"48",x"c0",x"e9",x"c1"),
  1406 => (x"41",x"20",x"49",x"6e"),
  1407 => (x"51",x"10",x"41",x"20"),
  1408 => (x"48",x"66",x"c4",x"c1"),
  1409 => (x"78",x"f3",x"d0",x"c1"),
  1410 => (x"81",x"c7",x"49",x"6a"),
  1411 => (x"c4",x"c1",x"51",x"74"),
  1412 => (x"81",x"c8",x"49",x"66"),
  1413 => (x"a6",x"d8",x"51",x"c1"),
  1414 => (x"c1",x"78",x"c2",x"48"),
  1415 => (x"c9",x"49",x"66",x"c4"),
  1416 => (x"c1",x"51",x"c0",x"81"),
  1417 => (x"ca",x"49",x"66",x"c4"),
  1418 => (x"c1",x"51",x"c0",x"81"),
  1419 => (x"6a",x"1e",x"d8",x"1e"),
  1420 => (x"ff",x"81",x"c8",x"49"),
  1421 => (x"c8",x"87",x"fa",x"df"),
  1422 => (x"66",x"c8",x"c1",x"86"),
  1423 => (x"01",x"a8",x"c0",x"48"),
  1424 => (x"a6",x"d0",x"87",x"c7"),
  1425 => (x"cf",x"78",x"c1",x"48"),
  1426 => (x"66",x"c8",x"c1",x"87"),
  1427 => (x"d8",x"88",x"c1",x"48"),
  1428 => (x"87",x"c4",x"58",x"a6"),
  1429 => (x"87",x"c5",x"df",x"ff"),
  1430 => (x"cd",x"02",x"9c",x"74"),
  1431 => (x"66",x"d0",x"87",x"da"),
  1432 => (x"66",x"cc",x"c1",x"48"),
  1433 => (x"cf",x"cd",x"03",x"a8"),
  1434 => (x"48",x"a6",x"c8",x"87"),
  1435 => (x"ff",x"7e",x"78",x"c0"),
  1436 => (x"70",x"87",x"c2",x"de"),
  1437 => (x"ac",x"d0",x"c1",x"4c"),
  1438 => (x"87",x"e7",x"c2",x"05"),
  1439 => (x"6e",x"48",x"a6",x"c4"),
  1440 => (x"87",x"d8",x"e0",x"78"),
  1441 => (x"cc",x"48",x"7e",x"70"),
  1442 => (x"c5",x"06",x"a8",x"66"),
  1443 => (x"48",x"a6",x"cc",x"87"),
  1444 => (x"dd",x"ff",x"78",x"6e"),
  1445 => (x"4c",x"70",x"87",x"df"),
  1446 => (x"05",x"ac",x"ec",x"c0"),
  1447 => (x"d0",x"87",x"ee",x"c1"),
  1448 => (x"91",x"cc",x"49",x"66"),
  1449 => (x"81",x"66",x"c4",x"c1"),
  1450 => (x"6a",x"4a",x"a1",x"c4"),
  1451 => (x"4a",x"a1",x"c8",x"4d"),
  1452 => (x"d1",x"c1",x"52",x"6e"),
  1453 => (x"dc",x"ff",x"79",x"f9"),
  1454 => (x"4c",x"70",x"87",x"fb"),
  1455 => (x"87",x"d9",x"02",x"9c"),
  1456 => (x"02",x"ac",x"fb",x"c0"),
  1457 => (x"55",x"74",x"87",x"d3"),
  1458 => (x"87",x"e9",x"dc",x"ff"),
  1459 => (x"02",x"9c",x"4c",x"70"),
  1460 => (x"fb",x"c0",x"87",x"c7"),
  1461 => (x"ed",x"ff",x"05",x"ac"),
  1462 => (x"55",x"e0",x"c0",x"87"),
  1463 => (x"c0",x"55",x"c1",x"c2"),
  1464 => (x"e0",x"c0",x"7d",x"97"),
  1465 => (x"66",x"c4",x"48",x"66"),
  1466 => (x"87",x"db",x"05",x"a8"),
  1467 => (x"d4",x"48",x"66",x"d0"),
  1468 => (x"ca",x"04",x"a8",x"66"),
  1469 => (x"48",x"66",x"d0",x"87"),
  1470 => (x"a6",x"d4",x"80",x"c1"),
  1471 => (x"d4",x"87",x"c8",x"58"),
  1472 => (x"88",x"c1",x"48",x"66"),
  1473 => (x"ff",x"58",x"a6",x"d8"),
  1474 => (x"70",x"87",x"ea",x"db"),
  1475 => (x"ac",x"d0",x"c1",x"4c"),
  1476 => (x"dc",x"87",x"c9",x"05"),
  1477 => (x"80",x"c1",x"48",x"66"),
  1478 => (x"58",x"a6",x"e0",x"c0"),
  1479 => (x"02",x"ac",x"d0",x"c1"),
  1480 => (x"6e",x"87",x"d9",x"fd"),
  1481 => (x"66",x"e0",x"c0",x"48"),
  1482 => (x"eb",x"c9",x"05",x"a8"),
  1483 => (x"a6",x"e4",x"c0",x"87"),
  1484 => (x"74",x"78",x"c0",x"48"),
  1485 => (x"88",x"fb",x"c0",x"48"),
  1486 => (x"70",x"58",x"a6",x"c8"),
  1487 => (x"dd",x"c9",x"02",x"98"),
  1488 => (x"88",x"cb",x"48",x"87"),
  1489 => (x"70",x"58",x"a6",x"c8"),
  1490 => (x"cf",x"c1",x"02",x"98"),
  1491 => (x"88",x"c9",x"48",x"87"),
  1492 => (x"70",x"58",x"a6",x"c8"),
  1493 => (x"ff",x"c3",x"02",x"98"),
  1494 => (x"88",x"c4",x"48",x"87"),
  1495 => (x"70",x"58",x"a6",x"c8"),
  1496 => (x"87",x"cf",x"02",x"98"),
  1497 => (x"c8",x"88",x"c1",x"48"),
  1498 => (x"98",x"70",x"58",x"a6"),
  1499 => (x"87",x"e8",x"c3",x"02"),
  1500 => (x"c8",x"87",x"dc",x"c8"),
  1501 => (x"f0",x"c0",x"48",x"a6"),
  1502 => (x"f8",x"d9",x"ff",x"78"),
  1503 => (x"c0",x"4c",x"70",x"87"),
  1504 => (x"c0",x"02",x"ac",x"ec"),
  1505 => (x"a6",x"cc",x"87",x"c3"),
  1506 => (x"ac",x"ec",x"c0",x"5c"),
  1507 => (x"ff",x"87",x"cd",x"02"),
  1508 => (x"70",x"87",x"e2",x"d9"),
  1509 => (x"ac",x"ec",x"c0",x"4c"),
  1510 => (x"87",x"f3",x"ff",x"05"),
  1511 => (x"02",x"ac",x"ec",x"c0"),
  1512 => (x"ff",x"87",x"c4",x"c0"),
  1513 => (x"c0",x"87",x"ce",x"d9"),
  1514 => (x"d8",x"1e",x"ca",x"1e"),
  1515 => (x"91",x"cc",x"49",x"66"),
  1516 => (x"48",x"66",x"cc",x"c1"),
  1517 => (x"a6",x"cc",x"80",x"71"),
  1518 => (x"48",x"66",x"c8",x"58"),
  1519 => (x"a6",x"d0",x"80",x"c4"),
  1520 => (x"bf",x"66",x"cc",x"58"),
  1521 => (x"e8",x"d9",x"ff",x"49"),
  1522 => (x"de",x"1e",x"c1",x"87"),
  1523 => (x"bf",x"66",x"d4",x"1e"),
  1524 => (x"dc",x"d9",x"ff",x"49"),
  1525 => (x"70",x"86",x"d0",x"87"),
  1526 => (x"08",x"c0",x"48",x"49"),
  1527 => (x"a6",x"ec",x"c0",x"88"),
  1528 => (x"06",x"a8",x"c0",x"58"),
  1529 => (x"c0",x"87",x"ee",x"c0"),
  1530 => (x"dd",x"48",x"66",x"e8"),
  1531 => (x"e4",x"c0",x"03",x"a8"),
  1532 => (x"bf",x"66",x"c4",x"87"),
  1533 => (x"66",x"e8",x"c0",x"49"),
  1534 => (x"51",x"e0",x"c0",x"81"),
  1535 => (x"49",x"66",x"e8",x"c0"),
  1536 => (x"66",x"c4",x"81",x"c1"),
  1537 => (x"c1",x"c2",x"81",x"bf"),
  1538 => (x"66",x"e8",x"c0",x"51"),
  1539 => (x"c4",x"81",x"c2",x"49"),
  1540 => (x"c0",x"81",x"bf",x"66"),
  1541 => (x"c1",x"48",x"6e",x"51"),
  1542 => (x"6e",x"78",x"f3",x"d0"),
  1543 => (x"d8",x"81",x"c8",x"49"),
  1544 => (x"49",x"6e",x"51",x"66"),
  1545 => (x"66",x"dc",x"81",x"c9"),
  1546 => (x"ca",x"49",x"6e",x"51"),
  1547 => (x"51",x"66",x"c8",x"81"),
  1548 => (x"c1",x"48",x"66",x"d8"),
  1549 => (x"58",x"a6",x"dc",x"80"),
  1550 => (x"d4",x"48",x"66",x"d0"),
  1551 => (x"c0",x"04",x"a8",x"66"),
  1552 => (x"66",x"d0",x"87",x"cb"),
  1553 => (x"d4",x"80",x"c1",x"48"),
  1554 => (x"d1",x"c5",x"58",x"a6"),
  1555 => (x"48",x"66",x"d4",x"87"),
  1556 => (x"a6",x"d8",x"88",x"c1"),
  1557 => (x"87",x"c6",x"c5",x"58"),
  1558 => (x"87",x"c0",x"d9",x"ff"),
  1559 => (x"58",x"a6",x"ec",x"c0"),
  1560 => (x"87",x"f8",x"d8",x"ff"),
  1561 => (x"58",x"a6",x"f0",x"c0"),
  1562 => (x"05",x"a8",x"ec",x"c0"),
  1563 => (x"a6",x"87",x"c9",x"c0"),
  1564 => (x"66",x"e8",x"c0",x"48"),
  1565 => (x"87",x"c4",x"c0",x"78"),
  1566 => (x"87",x"f9",x"d5",x"ff"),
  1567 => (x"cc",x"49",x"66",x"d0"),
  1568 => (x"66",x"c4",x"c1",x"91"),
  1569 => (x"c8",x"80",x"71",x"48"),
  1570 => (x"66",x"c4",x"58",x"a6"),
  1571 => (x"c4",x"82",x"c8",x"4a"),
  1572 => (x"81",x"ca",x"49",x"66"),
  1573 => (x"51",x"66",x"e8",x"c0"),
  1574 => (x"49",x"66",x"ec",x"c0"),
  1575 => (x"e8",x"c0",x"81",x"c1"),
  1576 => (x"48",x"c1",x"89",x"66"),
  1577 => (x"49",x"70",x"30",x"71"),
  1578 => (x"97",x"71",x"89",x"c1"),
  1579 => (x"c0",x"ee",x"c2",x"7a"),
  1580 => (x"e8",x"c0",x"49",x"bf"),
  1581 => (x"6a",x"97",x"29",x"66"),
  1582 => (x"98",x"71",x"48",x"4a"),
  1583 => (x"58",x"a6",x"f4",x"c0"),
  1584 => (x"c4",x"48",x"66",x"c4"),
  1585 => (x"58",x"a6",x"cc",x"80"),
  1586 => (x"4d",x"bf",x"66",x"c8"),
  1587 => (x"48",x"66",x"e0",x"c0"),
  1588 => (x"c0",x"02",x"a8",x"6e"),
  1589 => (x"7e",x"c0",x"87",x"c5"),
  1590 => (x"c1",x"87",x"c2",x"c0"),
  1591 => (x"c0",x"1e",x"6e",x"7e"),
  1592 => (x"49",x"75",x"1e",x"e0"),
  1593 => (x"87",x"c9",x"d5",x"ff"),
  1594 => (x"4c",x"70",x"86",x"c8"),
  1595 => (x"06",x"ac",x"b7",x"c0"),
  1596 => (x"74",x"87",x"d4",x"c1"),
  1597 => (x"bf",x"66",x"c8",x"85"),
  1598 => (x"81",x"e0",x"c0",x"49"),
  1599 => (x"c1",x"4b",x"89",x"75"),
  1600 => (x"71",x"4a",x"cc",x"e9"),
  1601 => (x"87",x"dc",x"e0",x"fe"),
  1602 => (x"7e",x"75",x"85",x"c2"),
  1603 => (x"48",x"66",x"e4",x"c0"),
  1604 => (x"e8",x"c0",x"80",x"c1"),
  1605 => (x"f0",x"c0",x"58",x"a6"),
  1606 => (x"81",x"c1",x"49",x"66"),
  1607 => (x"c0",x"02",x"a9",x"70"),
  1608 => (x"4d",x"c0",x"87",x"c5"),
  1609 => (x"c1",x"87",x"c2",x"c0"),
  1610 => (x"cc",x"1e",x"75",x"4d"),
  1611 => (x"c0",x"49",x"bf",x"66"),
  1612 => (x"66",x"c4",x"81",x"e0"),
  1613 => (x"c8",x"1e",x"71",x"89"),
  1614 => (x"d3",x"ff",x"49",x"66"),
  1615 => (x"86",x"c8",x"87",x"f3"),
  1616 => (x"01",x"a8",x"b7",x"c0"),
  1617 => (x"c0",x"87",x"c5",x"ff"),
  1618 => (x"c0",x"02",x"66",x"e4"),
  1619 => (x"66",x"c4",x"87",x"d3"),
  1620 => (x"c0",x"81",x"c9",x"49"),
  1621 => (x"c4",x"51",x"66",x"e4"),
  1622 => (x"d3",x"c1",x"48",x"66"),
  1623 => (x"ce",x"c0",x"78",x"c7"),
  1624 => (x"49",x"66",x"c4",x"87"),
  1625 => (x"51",x"c2",x"81",x"c9"),
  1626 => (x"c1",x"48",x"66",x"c4"),
  1627 => (x"d0",x"78",x"c5",x"d5"),
  1628 => (x"66",x"d4",x"48",x"66"),
  1629 => (x"cb",x"c0",x"04",x"a8"),
  1630 => (x"48",x"66",x"d0",x"87"),
  1631 => (x"a6",x"d4",x"80",x"c1"),
  1632 => (x"87",x"da",x"c0",x"58"),
  1633 => (x"c1",x"48",x"66",x"d4"),
  1634 => (x"58",x"a6",x"d8",x"88"),
  1635 => (x"ff",x"87",x"cf",x"c0"),
  1636 => (x"70",x"87",x"ca",x"d2"),
  1637 => (x"87",x"c6",x"c0",x"4c"),
  1638 => (x"87",x"c1",x"d2",x"ff"),
  1639 => (x"66",x"dc",x"4c",x"70"),
  1640 => (x"c0",x"80",x"c1",x"48"),
  1641 => (x"74",x"58",x"a6",x"e0"),
  1642 => (x"cb",x"c0",x"02",x"9c"),
  1643 => (x"48",x"66",x"d0",x"87"),
  1644 => (x"a8",x"66",x"cc",x"c1"),
  1645 => (x"87",x"f1",x"f2",x"04"),
  1646 => (x"c7",x"48",x"66",x"d0"),
  1647 => (x"e1",x"c0",x"03",x"a8"),
  1648 => (x"4c",x"66",x"d0",x"87"),
  1649 => (x"48",x"e4",x"ee",x"c2"),
  1650 => (x"49",x"74",x"78",x"c0"),
  1651 => (x"c4",x"c1",x"91",x"cc"),
  1652 => (x"a1",x"c4",x"81",x"66"),
  1653 => (x"c0",x"4a",x"6a",x"4a"),
  1654 => (x"84",x"c1",x"79",x"52"),
  1655 => (x"ff",x"04",x"ac",x"c7"),
  1656 => (x"e0",x"c0",x"87",x"e2"),
  1657 => (x"e2",x"c0",x"02",x"66"),
  1658 => (x"66",x"c4",x"c1",x"87"),
  1659 => (x"81",x"d4",x"c1",x"49"),
  1660 => (x"4a",x"66",x"c4",x"c1"),
  1661 => (x"c0",x"82",x"dc",x"c1"),
  1662 => (x"f9",x"d1",x"c1",x"52"),
  1663 => (x"66",x"c4",x"c1",x"79"),
  1664 => (x"81",x"d8",x"c1",x"49"),
  1665 => (x"79",x"d0",x"e9",x"c1"),
  1666 => (x"c1",x"87",x"d6",x"c0"),
  1667 => (x"c1",x"49",x"66",x"c4"),
  1668 => (x"c4",x"c1",x"81",x"d4"),
  1669 => (x"d8",x"c1",x"4a",x"66"),
  1670 => (x"d8",x"e9",x"c1",x"82"),
  1671 => (x"f0",x"d1",x"c1",x"7a"),
  1672 => (x"d7",x"d5",x"c1",x"79"),
  1673 => (x"66",x"c4",x"c1",x"4a"),
  1674 => (x"81",x"e0",x"c1",x"49"),
  1675 => (x"cf",x"ff",x"79",x"72"),
  1676 => (x"66",x"cc",x"87",x"e2"),
  1677 => (x"8e",x"cc",x"ff",x"48"),
  1678 => (x"4c",x"26",x"4d",x"26"),
  1679 => (x"4f",x"26",x"4b",x"26"),
  1680 => (x"64",x"61",x"6f",x"4c"),
  1681 => (x"20",x"2e",x"2a",x"20"),
  1682 => (x"00",x"00",x"00",x"00"),
  1683 => (x"00",x"00",x"20",x"3a"),
  1684 => (x"61",x"42",x"20",x"80"),
  1685 => (x"00",x"00",x"6b",x"63"),
  1686 => (x"78",x"45",x"20",x"80"),
  1687 => (x"1e",x"00",x"74",x"69"),
  1688 => (x"ee",x"c2",x"1e",x"c7"),
  1689 => (x"c1",x"1e",x"bf",x"e0"),
  1690 => (x"c2",x"1e",x"f0",x"ec"),
  1691 => (x"bf",x"97",x"c4",x"ee"),
  1692 => (x"87",x"f5",x"ec",x"49"),
  1693 => (x"49",x"f0",x"ec",x"c1"),
  1694 => (x"87",x"da",x"e1",x"c0"),
  1695 => (x"4f",x"26",x"8e",x"f4"),
  1696 => (x"c8",x"1e",x"73",x"1e"),
  1697 => (x"ee",x"c2",x"87",x"c3"),
  1698 => (x"50",x"c0",x"48",x"ec"),
  1699 => (x"48",x"c8",x"ee",x"c1"),
  1700 => (x"78",x"d0",x"ec",x"c1"),
  1701 => (x"49",x"a0",x"e8",x"fe"),
  1702 => (x"87",x"fa",x"e0",x"c0"),
  1703 => (x"e7",x"df",x"49",x"c7"),
  1704 => (x"c0",x"49",x"c1",x"87"),
  1705 => (x"ff",x"87",x"c2",x"e1"),
  1706 => (x"ff",x"c3",x"48",x"d4"),
  1707 => (x"db",x"e3",x"fe",x"78"),
  1708 => (x"02",x"98",x"70",x"87"),
  1709 => (x"ed",x"fe",x"87",x"cd"),
  1710 => (x"98",x"70",x"87",x"d7"),
  1711 => (x"c1",x"87",x"c4",x"02"),
  1712 => (x"c0",x"87",x"c2",x"4a"),
  1713 => (x"02",x"9a",x"72",x"4a"),
  1714 => (x"ec",x"c1",x"87",x"c8"),
  1715 => (x"d7",x"fe",x"49",x"dc"),
  1716 => (x"ee",x"c2",x"87",x"d5"),
  1717 => (x"78",x"c0",x"48",x"e0"),
  1718 => (x"48",x"c4",x"ee",x"c2"),
  1719 => (x"fd",x"49",x"50",x"c0"),
  1720 => (x"f4",x"c0",x"87",x"fd"),
  1721 => (x"4b",x"70",x"87",x"da"),
  1722 => (x"87",x"cb",x"02",x"9b"),
  1723 => (x"5b",x"cc",x"ee",x"c1"),
  1724 => (x"d3",x"de",x"49",x"c7"),
  1725 => (x"c0",x"87",x"c5",x"87"),
  1726 => (x"87",x"ed",x"df",x"49"),
  1727 => (x"c0",x"87",x"c4",x"c3"),
  1728 => (x"c0",x"87",x"ce",x"e1"),
  1729 => (x"ff",x"87",x"e2",x"ee"),
  1730 => (x"4b",x"26",x"87",x"f5"),
  1731 => (x"00",x"00",x"4f",x"26"),
  1732 => (x"74",x"6f",x"6f",x"42"),
  1733 => (x"2e",x"67",x"6e",x"69"),
  1734 => (x"00",x"00",x"2e",x"2e"),
  1735 => (x"4f",x"20",x"44",x"53"),
  1736 => (x"00",x"00",x"00",x"4b"),
  1737 => (x"00",x"00",x"00",x"00"),
  1738 => (x"00",x"00",x"00",x"00"),
  1739 => (x"00",x"00",x"00",x"01"),
  1740 => (x"00",x"00",x"11",x"5e"),
  1741 => (x"00",x"00",x"2b",x"b8"),
  1742 => (x"00",x"00",x"00",x"00"),
  1743 => (x"00",x"00",x"11",x"5e"),
  1744 => (x"00",x"00",x"2b",x"d6"),
  1745 => (x"00",x"00",x"00",x"00"),
  1746 => (x"00",x"00",x"11",x"5e"),
  1747 => (x"00",x"00",x"2b",x"f4"),
  1748 => (x"00",x"00",x"00",x"00"),
  1749 => (x"00",x"00",x"11",x"5e"),
  1750 => (x"00",x"00",x"2c",x"12"),
  1751 => (x"00",x"00",x"00",x"00"),
  1752 => (x"00",x"00",x"11",x"5e"),
  1753 => (x"00",x"00",x"2c",x"30"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"00",x"11",x"5e"),
  1756 => (x"00",x"00",x"2c",x"4e"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"11",x"5e"),
  1759 => (x"00",x"00",x"2c",x"6c"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"14",x"79"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"12",x"13"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"db",x"86",x"fc",x"1e"),
  1768 => (x"fc",x"7e",x"70",x"87"),
  1769 => (x"1e",x"4f",x"26",x"8e"),
  1770 => (x"c0",x"48",x"f0",x"fe"),
  1771 => (x"79",x"09",x"cd",x"78"),
  1772 => (x"1e",x"4f",x"26",x"09"),
  1773 => (x"49",x"dc",x"ee",x"c1"),
  1774 => (x"4f",x"26",x"87",x"ed"),
  1775 => (x"bf",x"f0",x"fe",x"1e"),
  1776 => (x"1e",x"4f",x"26",x"48"),
  1777 => (x"c1",x"48",x"f0",x"fe"),
  1778 => (x"1e",x"4f",x"26",x"78"),
  1779 => (x"c0",x"48",x"f0",x"fe"),
  1780 => (x"1e",x"4f",x"26",x"78"),
  1781 => (x"52",x"c0",x"4a",x"71"),
  1782 => (x"0e",x"4f",x"26",x"51"),
  1783 => (x"5d",x"5c",x"5b",x"5e"),
  1784 => (x"71",x"86",x"f4",x"0e"),
  1785 => (x"7e",x"6d",x"97",x"4d"),
  1786 => (x"97",x"4c",x"a5",x"c1"),
  1787 => (x"a6",x"c8",x"48",x"6c"),
  1788 => (x"c4",x"48",x"6e",x"58"),
  1789 => (x"c5",x"05",x"a8",x"66"),
  1790 => (x"c0",x"48",x"ff",x"87"),
  1791 => (x"ca",x"ff",x"87",x"e6"),
  1792 => (x"49",x"a5",x"c2",x"87"),
  1793 => (x"71",x"4b",x"6c",x"97"),
  1794 => (x"6b",x"97",x"4b",x"a3"),
  1795 => (x"7e",x"6c",x"97",x"4b"),
  1796 => (x"80",x"c1",x"48",x"6e"),
  1797 => (x"c7",x"58",x"a6",x"c8"),
  1798 => (x"58",x"a6",x"cc",x"98"),
  1799 => (x"fe",x"7c",x"97",x"70"),
  1800 => (x"48",x"73",x"87",x"e1"),
  1801 => (x"4d",x"26",x"8e",x"f4"),
  1802 => (x"4b",x"26",x"4c",x"26"),
  1803 => (x"5e",x"0e",x"4f",x"26"),
  1804 => (x"f4",x"0e",x"5c",x"5b"),
  1805 => (x"d8",x"4c",x"71",x"86"),
  1806 => (x"ff",x"c3",x"4a",x"66"),
  1807 => (x"4b",x"a4",x"c2",x"9a"),
  1808 => (x"73",x"49",x"6c",x"97"),
  1809 => (x"51",x"72",x"49",x"a1"),
  1810 => (x"6e",x"7e",x"6c",x"97"),
  1811 => (x"c8",x"80",x"c1",x"48"),
  1812 => (x"98",x"c7",x"58",x"a6"),
  1813 => (x"70",x"58",x"a6",x"cc"),
  1814 => (x"26",x"8e",x"f4",x"54"),
  1815 => (x"26",x"4b",x"26",x"4c"),
  1816 => (x"86",x"fc",x"1e",x"4f"),
  1817 => (x"e0",x"87",x"e4",x"fd"),
  1818 => (x"c0",x"49",x"4a",x"bf"),
  1819 => (x"02",x"99",x"c0",x"e0"),
  1820 => (x"1e",x"72",x"87",x"cb"),
  1821 => (x"49",x"cc",x"f2",x"c2"),
  1822 => (x"c4",x"87",x"f3",x"fe"),
  1823 => (x"87",x"fc",x"fc",x"86"),
  1824 => (x"fe",x"fc",x"7e",x"70"),
  1825 => (x"26",x"8e",x"fc",x"87"),
  1826 => (x"f2",x"c2",x"1e",x"4f"),
  1827 => (x"c2",x"fd",x"49",x"cc"),
  1828 => (x"e1",x"f1",x"c1",x"87"),
  1829 => (x"87",x"cf",x"fc",x"49"),
  1830 => (x"26",x"87",x"f1",x"c2"),
  1831 => (x"1e",x"73",x"1e",x"4f"),
  1832 => (x"49",x"cc",x"f2",x"c2"),
  1833 => (x"70",x"87",x"f4",x"fc"),
  1834 => (x"aa",x"b7",x"c0",x"4a"),
  1835 => (x"87",x"cc",x"c2",x"04"),
  1836 => (x"05",x"aa",x"f0",x"c3"),
  1837 => (x"f5",x"c1",x"87",x"c9"),
  1838 => (x"78",x"c1",x"48",x"c4"),
  1839 => (x"c3",x"87",x"ed",x"c1"),
  1840 => (x"c9",x"05",x"aa",x"e0"),
  1841 => (x"c8",x"f5",x"c1",x"87"),
  1842 => (x"c1",x"78",x"c1",x"48"),
  1843 => (x"f5",x"c1",x"87",x"de"),
  1844 => (x"c6",x"02",x"bf",x"c8"),
  1845 => (x"a2",x"c0",x"c2",x"87"),
  1846 => (x"72",x"87",x"c2",x"4b"),
  1847 => (x"c4",x"f5",x"c1",x"4b"),
  1848 => (x"e0",x"c0",x"02",x"bf"),
  1849 => (x"c4",x"49",x"73",x"87"),
  1850 => (x"c1",x"91",x"29",x"b7"),
  1851 => (x"73",x"81",x"e0",x"f6"),
  1852 => (x"c2",x"9a",x"cf",x"4a"),
  1853 => (x"72",x"48",x"c1",x"92"),
  1854 => (x"ff",x"4a",x"70",x"30"),
  1855 => (x"69",x"48",x"72",x"ba"),
  1856 => (x"db",x"79",x"70",x"98"),
  1857 => (x"c4",x"49",x"73",x"87"),
  1858 => (x"c1",x"91",x"29",x"b7"),
  1859 => (x"73",x"81",x"e0",x"f6"),
  1860 => (x"c2",x"9a",x"cf",x"4a"),
  1861 => (x"72",x"48",x"c3",x"92"),
  1862 => (x"48",x"4a",x"70",x"30"),
  1863 => (x"79",x"70",x"b0",x"69"),
  1864 => (x"48",x"c8",x"f5",x"c1"),
  1865 => (x"f5",x"c1",x"78",x"c0"),
  1866 => (x"78",x"c0",x"48",x"c4"),
  1867 => (x"49",x"cc",x"f2",x"c2"),
  1868 => (x"70",x"87",x"e8",x"fa"),
  1869 => (x"aa",x"b7",x"c0",x"4a"),
  1870 => (x"87",x"f4",x"fd",x"03"),
  1871 => (x"4b",x"26",x"48",x"c0"),
  1872 => (x"00",x"00",x"4f",x"26"),
  1873 => (x"00",x"00",x"00",x"00"),
  1874 => (x"00",x"00",x"00",x"00"),
  1875 => (x"72",x"4a",x"c0",x"1e"),
  1876 => (x"c1",x"91",x"c4",x"49"),
  1877 => (x"c0",x"81",x"e0",x"f6"),
  1878 => (x"d0",x"82",x"c1",x"79"),
  1879 => (x"ee",x"04",x"aa",x"b7"),
  1880 => (x"0e",x"4f",x"26",x"87"),
  1881 => (x"5d",x"5c",x"5b",x"5e"),
  1882 => (x"f9",x"4d",x"71",x"0e"),
  1883 => (x"4a",x"75",x"87",x"dd"),
  1884 => (x"92",x"2a",x"b7",x"c4"),
  1885 => (x"82",x"e0",x"f6",x"c1"),
  1886 => (x"9c",x"cf",x"4c",x"75"),
  1887 => (x"49",x"6a",x"94",x"c2"),
  1888 => (x"c3",x"2b",x"74",x"4b"),
  1889 => (x"74",x"48",x"c2",x"9b"),
  1890 => (x"ff",x"4c",x"70",x"30"),
  1891 => (x"71",x"48",x"74",x"bc"),
  1892 => (x"f8",x"7a",x"70",x"98"),
  1893 => (x"48",x"73",x"87",x"ed"),
  1894 => (x"4c",x"26",x"4d",x"26"),
  1895 => (x"4f",x"26",x"4b",x"26"),
  1896 => (x"00",x"00",x"00",x"00"),
  1897 => (x"00",x"00",x"00",x"00"),
  1898 => (x"00",x"00",x"00",x"00"),
  1899 => (x"00",x"00",x"00",x"00"),
  1900 => (x"00",x"00",x"00",x"00"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"00",x"00",x"00",x"00"),
  1904 => (x"00",x"00",x"00",x"00"),
  1905 => (x"00",x"00",x"00",x"00"),
  1906 => (x"00",x"00",x"00",x"00"),
  1907 => (x"00",x"00",x"00",x"00"),
  1908 => (x"00",x"00",x"00",x"00"),
  1909 => (x"00",x"00",x"00",x"00"),
  1910 => (x"00",x"00",x"00",x"00"),
  1911 => (x"00",x"00",x"00",x"00"),
  1912 => (x"48",x"d0",x"ff",x"1e"),
  1913 => (x"71",x"78",x"e1",x"c8"),
  1914 => (x"08",x"d4",x"ff",x"48"),
  1915 => (x"1e",x"4f",x"26",x"78"),
  1916 => (x"c8",x"48",x"d0",x"ff"),
  1917 => (x"48",x"71",x"78",x"e1"),
  1918 => (x"78",x"08",x"d4",x"ff"),
  1919 => (x"ff",x"48",x"66",x"c4"),
  1920 => (x"26",x"78",x"08",x"d4"),
  1921 => (x"4a",x"71",x"1e",x"4f"),
  1922 => (x"1e",x"49",x"66",x"c4"),
  1923 => (x"de",x"ff",x"49",x"72"),
  1924 => (x"48",x"d0",x"ff",x"87"),
  1925 => (x"fc",x"78",x"e0",x"c0"),
  1926 => (x"1e",x"4f",x"26",x"8e"),
  1927 => (x"4b",x"71",x"1e",x"73"),
  1928 => (x"1e",x"49",x"66",x"c8"),
  1929 => (x"e0",x"c1",x"4a",x"73"),
  1930 => (x"d8",x"ff",x"49",x"a2"),
  1931 => (x"26",x"8e",x"fc",x"87"),
  1932 => (x"1e",x"4f",x"26",x"4b"),
  1933 => (x"c8",x"48",x"d0",x"ff"),
  1934 => (x"48",x"71",x"78",x"c9"),
  1935 => (x"78",x"08",x"d4",x"ff"),
  1936 => (x"71",x"1e",x"4f",x"26"),
  1937 => (x"87",x"eb",x"49",x"4a"),
  1938 => (x"c8",x"48",x"d0",x"ff"),
  1939 => (x"1e",x"4f",x"26",x"78"),
  1940 => (x"4b",x"71",x"1e",x"73"),
  1941 => (x"bf",x"e4",x"f2",x"c2"),
  1942 => (x"c2",x"87",x"c3",x"02"),
  1943 => (x"d0",x"ff",x"87",x"eb"),
  1944 => (x"78",x"c9",x"c8",x"48"),
  1945 => (x"e0",x"c0",x"48",x"73"),
  1946 => (x"08",x"d4",x"ff",x"b0"),
  1947 => (x"d8",x"f2",x"c2",x"78"),
  1948 => (x"c8",x"78",x"c0",x"48"),
  1949 => (x"87",x"c5",x"02",x"66"),
  1950 => (x"c2",x"49",x"ff",x"c3"),
  1951 => (x"c2",x"49",x"c0",x"87"),
  1952 => (x"cc",x"59",x"e0",x"f2"),
  1953 => (x"87",x"c6",x"02",x"66"),
  1954 => (x"4a",x"d5",x"d5",x"c5"),
  1955 => (x"ff",x"cf",x"87",x"c4"),
  1956 => (x"f2",x"c2",x"4a",x"ff"),
  1957 => (x"f2",x"c2",x"5a",x"e4"),
  1958 => (x"78",x"c1",x"48",x"e4"),
  1959 => (x"4f",x"26",x"4b",x"26"),
  1960 => (x"5c",x"5b",x"5e",x"0e"),
  1961 => (x"4d",x"71",x"0e",x"5d"),
  1962 => (x"bf",x"e0",x"f2",x"c2"),
  1963 => (x"02",x"9d",x"75",x"4b"),
  1964 => (x"c8",x"49",x"87",x"cb"),
  1965 => (x"c8",x"f9",x"c1",x"91"),
  1966 => (x"c4",x"82",x"71",x"4a"),
  1967 => (x"c8",x"fd",x"c1",x"87"),
  1968 => (x"12",x"4c",x"c0",x"4a"),
  1969 => (x"c2",x"99",x"73",x"49"),
  1970 => (x"48",x"bf",x"dc",x"f2"),
  1971 => (x"d4",x"ff",x"b8",x"71"),
  1972 => (x"b7",x"c1",x"78",x"08"),
  1973 => (x"b7",x"c8",x"84",x"2b"),
  1974 => (x"87",x"e7",x"04",x"ac"),
  1975 => (x"bf",x"d8",x"f2",x"c2"),
  1976 => (x"c2",x"80",x"c8",x"48"),
  1977 => (x"26",x"58",x"dc",x"f2"),
  1978 => (x"26",x"4c",x"26",x"4d"),
  1979 => (x"1e",x"4f",x"26",x"4b"),
  1980 => (x"4b",x"71",x"1e",x"73"),
  1981 => (x"02",x"9a",x"4a",x"13"),
  1982 => (x"49",x"72",x"87",x"cb"),
  1983 => (x"13",x"87",x"e1",x"fe"),
  1984 => (x"f5",x"05",x"9a",x"4a"),
  1985 => (x"26",x"4b",x"26",x"87"),
  1986 => (x"f2",x"c2",x"1e",x"4f"),
  1987 => (x"c2",x"49",x"bf",x"d8"),
  1988 => (x"c1",x"48",x"d8",x"f2"),
  1989 => (x"c0",x"c4",x"78",x"a1"),
  1990 => (x"db",x"03",x"a9",x"b7"),
  1991 => (x"48",x"d4",x"ff",x"87"),
  1992 => (x"bf",x"dc",x"f2",x"c2"),
  1993 => (x"d8",x"f2",x"c2",x"78"),
  1994 => (x"f2",x"c2",x"49",x"bf"),
  1995 => (x"a1",x"c1",x"48",x"d8"),
  1996 => (x"b7",x"c0",x"c4",x"78"),
  1997 => (x"87",x"e5",x"04",x"a9"),
  1998 => (x"c8",x"48",x"d0",x"ff"),
  1999 => (x"e4",x"f2",x"c2",x"78"),
  2000 => (x"26",x"78",x"c0",x"48"),
  2001 => (x"00",x"00",x"00",x"4f"),
  2002 => (x"00",x"00",x"00",x"00"),
  2003 => (x"00",x"00",x"00",x"00"),
  2004 => (x"5f",x"00",x"00",x"00"),
  2005 => (x"00",x"00",x"00",x"5f"),
  2006 => (x"00",x"03",x"03",x"00"),
  2007 => (x"00",x"00",x"03",x"03"),
  2008 => (x"14",x"7f",x"7f",x"14"),
  2009 => (x"00",x"14",x"7f",x"7f"),
  2010 => (x"6b",x"2e",x"24",x"00"),
  2011 => (x"00",x"12",x"3a",x"6b"),
  2012 => (x"18",x"36",x"6a",x"4c"),
  2013 => (x"00",x"32",x"56",x"6c"),
  2014 => (x"59",x"4f",x"7e",x"30"),
  2015 => (x"40",x"68",x"3a",x"77"),
  2016 => (x"07",x"04",x"00",x"00"),
  2017 => (x"00",x"00",x"00",x"03"),
  2018 => (x"3e",x"1c",x"00",x"00"),
  2019 => (x"00",x"00",x"41",x"63"),
  2020 => (x"63",x"41",x"00",x"00"),
  2021 => (x"00",x"00",x"1c",x"3e"),
  2022 => (x"1c",x"3e",x"2a",x"08"),
  2023 => (x"08",x"2a",x"3e",x"1c"),
  2024 => (x"3e",x"08",x"08",x"00"),
  2025 => (x"00",x"08",x"08",x"3e"),
  2026 => (x"e0",x"80",x"00",x"00"),
  2027 => (x"00",x"00",x"00",x"60"),
  2028 => (x"08",x"08",x"08",x"00"),
  2029 => (x"00",x"08",x"08",x"08"),
  2030 => (x"60",x"00",x"00",x"00"),
  2031 => (x"00",x"00",x"00",x"60"),
  2032 => (x"18",x"30",x"60",x"40"),
  2033 => (x"01",x"03",x"06",x"0c"),
  2034 => (x"59",x"7f",x"3e",x"00"),
  2035 => (x"00",x"3e",x"7f",x"4d"),
  2036 => (x"7f",x"06",x"04",x"00"),
  2037 => (x"00",x"00",x"00",x"7f"),
  2038 => (x"71",x"63",x"42",x"00"),
  2039 => (x"00",x"46",x"4f",x"59"),
  2040 => (x"49",x"63",x"22",x"00"),
  2041 => (x"00",x"36",x"7f",x"49"),
  2042 => (x"13",x"16",x"1c",x"18"),
  2043 => (x"00",x"10",x"7f",x"7f"),
  2044 => (x"45",x"67",x"27",x"00"),
  2045 => (x"00",x"39",x"7d",x"45"),
  2046 => (x"4b",x"7e",x"3c",x"00"),
  2047 => (x"00",x"30",x"79",x"49"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

